localparam [63:0] WBL_ROM1 [0:63] = '{
    64'h55bbc9a1bacd0963,
    64'hd445fb36780c837c,
    64'hc753bc0025132c77,
    64'h000000002eec1a7b,
    64'h000000001c5f1bf2,
    64'h00000000a6976e6b,
    64'h00000000b4445a6f,
    64'h00000000c617a0c5,
    64'h00000000e8c45230,
    64'h00000000dda73b01,
    64'h00000000747ed667,
    64'h000000001f3db32b,
    64'h000000004b6429fe,
    64'h00000000bd5de3d7,
    64'h000000008b192fab,
    64'h000000008a738476,
    64'h00000000706053ca,
    64'h000000003e81d182,
    64'h00000000b54f00c9,
    64'h0000000066dced7d,
    64'h00000000482220fa,
    64'h00000000032afc59,
    64'h00000000f690b147,
    64'h000000000e885bf0,
    64'h0000000061466aad,
    64'h0000000035eecbd4,
    64'h0000000057b8bea2,
    64'h00000000b91439af,
    64'h0000000086de4a9c,
    64'h00000000c15e4ca4,
    64'h000000001d0b5872,
    64'h000000009edbcfc0,
    64'haa44365ee1e0d0b7,
    64'h2bba04c9f832effd,
    64'h38ac4300983aaa93,
    64'h00000000110afb26,
    64'h0000000069494336,
    64'h00000000d9064d3f,
    64'h000000008e2433f7,
    64'h00000000945c85cc,
    64'h000000009bc24534,
    64'h000000001ed3f9a5,
    64'h0000000087ac02e5,
    64'h00000000e9627ff1,
    64'h00000000ce915071,
    64'h0000000055953cd8,
    64'h0000000028e49f31,
    64'h00000000df79a815,
    64'h000000008ce75104,
    64'h00000000a1c8a3c7,
    64'h0000000089374023,
    64'h000000000d6d8fc3,
    64'h00000000bf8d9218,
    64'h00000000e6d59d96,
    64'h00000000424e3805,
    64'h0000000068a9f59a,
    64'h00000000416cbc07,
    64'h000000009956b612,
    64'h000000002df4da80,
    64'h000000000fea21e2,
    64'h00000000b06510eb,
    64'h00000000547aff27,
    64'h00000000bbaef3b2,
    64'h000000001608d275
};

localparam [63:0] WBL_ROM2 [0:63] = '{
    64'h33c3fccfbacd0963,
    64'hf396ed8e780c837c,
    64'hf297460025132c77,
    64'h000000002eec1a7b,
    64'h000000001c5f1bf2,
    64'h00000000a6976e6b,
    64'h00000000b4445a6f,
    64'h00000000c617a0c5,
    64'h00000000e8c45230,
    64'h00000000dda73b01,
    64'h00000000747ed667,
    64'h000000001f3db32b,
    64'h000000004b6429fe,
    64'h00000000bd5de3d7,
    64'h000000008b192fab,
    64'h000000008a738476,
    64'h00000000706053ca,
    64'h000000003e81d182,
    64'h00000000b54f00c9,
    64'h0000000066dced7d,
    64'h00000000482220fa,
    64'h00000000032afc59,
    64'h00000000f690b147,
    64'h000000000e885bf0,
    64'h0000000061466aad,
    64'h0000000035eecbd4,
    64'h0000000057b8bea2,
    64'h00000000b91439af,
    64'h0000000086de4a9c,
    64'h00000000c15e4ca4,
    64'h000000001d0b5872,
    64'h000000009edbcfc0,
    64'hcc3c0330e1e0d0b7,
    64'h0c691271f832effd,
    64'h0d68b900983aaa93,
    64'h00000000110afb26,
    64'h0000000069494336,
    64'h00000000d9064d3f,
    64'h000000008e2433f7,
    64'h00000000945c85cc,
    64'h000000009bc24534,
    64'h000000001ed3f9a5,
    64'h0000000087ac02e5,
    64'h00000000e9627ff1,
    64'h00000000ce915071,
    64'h0000000055953cd8,
    64'h0000000028e49f31,
    64'h00000000df79a815,
    64'h000000008ce75104,
    64'h00000000a1c8a3c7,
    64'h0000000089374023,
    64'h000000000d6d8fc3,
    64'h00000000bf8d9218,
    64'h00000000e6d59d96,
    64'h00000000424e3805,
    64'h0000000068a9f59a,
    64'h00000000416cbc07,
    64'h000000009956b612,
    64'h000000002df4da80,
    64'h000000000fea21e2,
    64'h00000000b06510eb,
    64'h00000000547aff27,
    64'h00000000bbaef3b2,
    64'h000000001608d275
};

localparam [63:0] WBL_ROM3 [0:63] = '{
    64'h0f0c5a1dbacd0963,
    64'h1bb6c706780c837c,
    64'h0706520025132c77,
    64'h000000002eec1a7b,
    64'h000000001c5f1bf2,
    64'h00000000a6976e6b,
    64'h00000000b4445a6f,
    64'h00000000c617a0c5,
    64'h00000000e8c45230,
    64'h00000000dda73b01,
    64'h00000000747ed667,
    64'h000000001f3db32b,
    64'h000000004b6429fe,
    64'h00000000bd5de3d7,
    64'h000000008b192fab,
    64'h000000008a738476,
    64'h00000000706053ca,
    64'h000000003e81d182,
    64'h00000000b54f00c9,
    64'h0000000066dced7d,
    64'h00000000482220fa,
    64'h00000000032afc59,
    64'h00000000f690b147,
    64'h000000000e885bf0,
    64'h0000000061466aad,
    64'h0000000035eecbd4,
    64'h0000000057b8bea2,
    64'h00000000b91439af,
    64'h0000000086de4a9c,
    64'h00000000c15e4ca4,
    64'h000000001d0b5872,
    64'h000000009edbcfc0,
    64'hf0f3a5e2e1e0d0b7,
    64'he44938f9f832effd,
    64'hf8f9ad00983aaa93,
    64'h00000000110afb26,
    64'h0000000069494336,
    64'h00000000d9064d3f,
    64'h000000008e2433f7,
    64'h00000000945c85cc,
    64'h000000009bc24534,
    64'h000000001ed3f9a5,
    64'h0000000087ac02e5,
    64'h00000000e9627ff1,
    64'h00000000ce915071,
    64'h0000000055953cd8,
    64'h0000000028e49f31,
    64'h00000000df79a815,
    64'h000000008ce75104,
    64'h00000000a1c8a3c7,
    64'h0000000089374023,
    64'h000000000d6d8fc3,
    64'h00000000bf8d9218,
    64'h00000000e6d59d96,
    64'h00000000424e3805,
    64'h0000000068a9f59a,
    64'h00000000416cbc07,
    64'h000000009956b612,
    64'h000000002df4da80,
    64'h000000000fea21e2,
    64'h00000000b06510eb,
    64'h00000000547aff27,
    64'h00000000bbaef3b2,
    64'h000000001608d275
};

localparam [63:0] WBL_ROM4 [0:63] = '{
    64'h00ff99e1bacd0963,
    64'h7e98b5c4780c837c,
    64'h05fbc90025132c77,
    64'h000000002eec1a7b,
    64'h000000001c5f1bf2,
    64'h00000000a6976e6b,
    64'h00000000b4445a6f,
    64'h00000000c617a0c5,
    64'h00000000e8c45230,
    64'h00000000dda73b01,
    64'h00000000747ed667,
    64'h000000001f3db32b,
    64'h000000004b6429fe,
    64'h00000000bd5de3d7,
    64'h000000008b192fab,
    64'h000000008a738476,
    64'h00000000706053ca,
    64'h000000003e81d182,
    64'h00000000b54f00c9,
    64'h0000000066dced7d,
    64'h00000000482220fa,
    64'h00000000032afc59,
    64'h00000000f690b147,
    64'h000000000e885bf0,
    64'h0000000061466aad,
    64'h0000000035eecbd4,
    64'h0000000057b8bea2,
    64'h00000000b91439af,
    64'h0000000086de4a9c,
    64'h00000000c15e4ca4,
    64'h000000001d0b5872,
    64'h000000009edbcfc0,
    64'hff00661ee1e0d0b7,
    64'h81674a3bf832effd,
    64'hfa043600983aaa93,
    64'h00000000110afb26,
    64'h0000000069494336,
    64'h00000000d9064d3f,
    64'h000000008e2433f7,
    64'h00000000945c85cc,
    64'h000000009bc24534,
    64'h000000001ed3f9a5,
    64'h0000000087ac02e5,
    64'h00000000e9627ff1,
    64'h00000000ce915071,
    64'h0000000055953cd8,
    64'h0000000028e49f31,
    64'h00000000df79a815,
    64'h000000008ce75104,
    64'h00000000a1c8a3c7,
    64'h0000000089374023,
    64'h000000000d6d8fc3,
    64'h00000000bf8d9218,
    64'h00000000e6d59d96,
    64'h00000000424e3805,
    64'h0000000068a9f59a,
    64'h00000000416cbc07,
    64'h000000009956b612,
    64'h000000002df4da80,
    64'h000000000fea21e2,
    64'h00000000b06510eb,
    64'h00000000547aff27,
    64'h00000000bbaef3b2,
    64'h000000001608d275
};

localparam [63:0] WBL_ROM5 [0:63] = '{
    64'h0055bbc9bacd0963,
    64'h5ee72c70780c837c,
    64'h3f662d0025132c77,
    64'h000000002eec1a7b,
    64'h000000001c5f1bf2,
    64'h00000000a6976e6b,
    64'h00000000b4445a6f,
    64'h00000000c617a0c5,
    64'h00000000e8c45230,
    64'h00000000dda73b01,
    64'h00000000747ed667,
    64'h000000001f3db32b,
    64'h000000004b6429fe,
    64'h00000000bd5de3d7,
    64'h000000008b192fab,
    64'h000000008a738476,
    64'h00000000706053ca,
    64'h000000003e81d182,
    64'h00000000b54f00c9,
    64'h0000000066dced7d,
    64'h00000000482220fa,
    64'h00000000032afc59,
    64'h00000000f690b147,
    64'h000000000e885bf0,
    64'h0000000061466aad,
    64'h0000000035eecbd4,
    64'h0000000057b8bea2,
    64'h00000000b91439af,
    64'h0000000086de4a9c,
    64'h00000000c15e4ca4,
    64'h000000001d0b5872,
    64'h000000009edbcfc0,
    64'hffaa4436e1e0d0b7,
    64'ha118d38ff832effd,
    64'hc099d200983aaa93,
    64'h00000000110afb26,
    64'h0000000069494336,
    64'h00000000d9064d3f,
    64'h000000008e2433f7,
    64'h00000000945c85cc,
    64'h000000009bc24534,
    64'h000000001ed3f9a5,
    64'h0000000087ac02e5,
    64'h00000000e9627ff1,
    64'h00000000ce915071,
    64'h0000000055953cd8,
    64'h0000000028e49f31,
    64'h00000000df79a815,
    64'h000000008ce75104,
    64'h00000000a1c8a3c7,
    64'h0000000089374023,
    64'h000000000d6d8fc3,
    64'h00000000bf8d9218,
    64'h00000000e6d59d96,
    64'h00000000424e3805,
    64'h0000000068a9f59a,
    64'h00000000416cbc07,
    64'h000000009956b612,
    64'h000000002df4da80,
    64'h000000000fea21e2,
    64'h00000000b06510eb,
    64'h00000000547aff27,
    64'h00000000bbaef3b2,
    64'h000000001608d275
};

localparam [63:0] WBL_ROM6 [0:63] = '{
    64'h00ff6678bacd0963,
    64'hca08a07f780c837c,
    64'h99b43a0025132c77,
    64'h000000002eec1a7b,
    64'h000000001c5f1bf2,
    64'h00000000a6976e6b,
    64'h00000000b4445a6f,
    64'h00000000c617a0c5,
    64'h00000000e8c45230,
    64'h00000000dda73b01,
    64'h00000000747ed667,
    64'h000000001f3db32b,
    64'h000000004b6429fe,
    64'h00000000bd5de3d7,
    64'h000000008b192fab,
    64'h000000008a738476,
    64'h00000000706053ca,
    64'h000000003e81d182,
    64'h00000000b54f00c9,
    64'h0000000066dced7d,
    64'h00000000482220fa,
    64'h00000000032afc59,
    64'h00000000f690b147,
    64'h000000000e885bf0,
    64'h0000000061466aad,
    64'h0000000035eecbd4,
    64'h0000000057b8bea2,
    64'h00000000b91439af,
    64'h0000000086de4a9c,
    64'h00000000c15e4ca4,
    64'h000000001d0b5872,
    64'h000000009edbcfc0,
    64'hff009987e1e0d0b7,
    64'h35f75f80f832effd,
    64'h664bc500983aaa93,
    64'h00000000110afb26,
    64'h0000000069494336,
    64'h00000000d9064d3f,
    64'h000000008e2433f7,
    64'h00000000945c85cc,
    64'h000000009bc24534,
    64'h000000001ed3f9a5,
    64'h0000000087ac02e5,
    64'h00000000e9627ff1,
    64'h00000000ce915071,
    64'h0000000055953cd8,
    64'h0000000028e49f31,
    64'h00000000df79a815,
    64'h000000008ce75104,
    64'h00000000a1c8a3c7,
    64'h0000000089374023,
    64'h000000000d6d8fc3,
    64'h00000000bf8d9218,
    64'h00000000e6d59d96,
    64'h00000000424e3805,
    64'h0000000068a9f59a,
    64'h00000000416cbc07,
    64'h000000009956b612,
    64'h000000002df4da80,
    64'h000000000fea21e2,
    64'h00000000b06510eb,
    64'h00000000547aff27,
    64'h00000000bbaef3b2,
    64'h000000001608d275
};

localparam [63:0] WBL_ROM7 [0:63] = '{
    64'h00aaddb1bacd0963,
    64'h6b763835780c837c,
    64'h6e272c0025132c77,
    64'h000000002eec1a7b,
    64'h000000001c5f1bf2,
    64'h00000000a6976e6b,
    64'h00000000b4445a6f,
    64'h00000000c617a0c5,
    64'h00000000e8c45230,
    64'h00000000dda73b01,
    64'h00000000747ed667,
    64'h000000001f3db32b,
    64'h000000004b6429fe,
    64'h00000000bd5de3d7,
    64'h000000008b192fab,
    64'h000000008a738476,
    64'h00000000706053ca,
    64'h000000003e81d182,
    64'h00000000b54f00c9,
    64'h0000000066dced7d,
    64'h00000000482220fa,
    64'h00000000032afc59,
    64'h00000000f690b147,
    64'h000000000e885bf0,
    64'h0000000061466aad,
    64'h0000000035eecbd4,
    64'h0000000057b8bea2,
    64'h00000000b91439af,
    64'h0000000086de4a9c,
    64'h00000000c15e4ca4,
    64'h000000001d0b5872,
    64'h000000009edbcfc0,
    64'hff55224ee1e0d0b7,
    64'h9489c7caf832effd,
    64'h91d8d300983aaa93,
    64'h00000000110afb26,
    64'h0000000069494336,
    64'h00000000d9064d3f,
    64'h000000008e2433f7,
    64'h00000000945c85cc,
    64'h000000009bc24534,
    64'h000000001ed3f9a5,
    64'h0000000087ac02e5,
    64'h00000000e9627ff1,
    64'h00000000ce915071,
    64'h0000000055953cd8,
    64'h0000000028e49f31,
    64'h00000000df79a815,
    64'h000000008ce75104,
    64'h00000000a1c8a3c7,
    64'h0000000089374023,
    64'h000000000d6d8fc3,
    64'h00000000bf8d9218,
    64'h00000000e6d59d96,
    64'h00000000424e3805,
    64'h0000000068a9f59a,
    64'h00000000416cbc07,
    64'h000000009956b612,
    64'h000000002df4da80,
    64'h000000000fea21e2,
    64'h00000000b06510eb,
    64'h00000000547aff27,
    64'h00000000bbaef3b2,
    64'h000000001608d275
};

localparam [63:0] WBL_ROM8 [0:63] = '{
    64'h00005511bacd0963,
    64'heb766d24780c837c,
    64'hd015ee0025132c77,
    64'h000000002eec1a7b,
    64'h000000001c5f1bf2,
    64'h00000000a6976e6b,
    64'h00000000b4445a6f,
    64'h00000000c617a0c5,
    64'h00000000e8c45230,
    64'h00000000dda73b01,
    64'h00000000747ed667,
    64'h000000001f3db32b,
    64'h000000004b6429fe,
    64'h00000000bd5de3d7,
    64'h000000008b192fab,
    64'h000000008a738476,
    64'h00000000706053ca,
    64'h000000003e81d182,
    64'h00000000b54f00c9,
    64'h0000000066dced7d,
    64'h00000000482220fa,
    64'h00000000032afc59,
    64'h00000000f690b147,
    64'h000000000e885bf0,
    64'h0000000061466aad,
    64'h0000000035eecbd4,
    64'h0000000057b8bea2,
    64'h00000000b91439af,
    64'h0000000086de4a9c,
    64'h00000000c15e4ca4,
    64'h000000001d0b5872,
    64'h000000009edbcfc0,
    64'hffffaaeee1e0d0b7,
    64'h148992dbf832effd,
    64'h2fea1100983aaa93,
    64'h00000000110afb26,
    64'h0000000069494336,
    64'h00000000d9064d3f,
    64'h000000008e2433f7,
    64'h00000000945c85cc,
    64'h000000009bc24534,
    64'h000000001ed3f9a5,
    64'h0000000087ac02e5,
    64'h00000000e9627ff1,
    64'h00000000ce915071,
    64'h0000000055953cd8,
    64'h0000000028e49f31,
    64'h00000000df79a815,
    64'h000000008ce75104,
    64'h00000000a1c8a3c7,
    64'h0000000089374023,
    64'h000000000d6d8fc3,
    64'h00000000bf8d9218,
    64'h00000000e6d59d96,
    64'h00000000424e3805,
    64'h0000000068a9f59a,
    64'h00000000416cbc07,
    64'h000000009956b612,
    64'h000000002df4da80,
    64'h000000000fea21e2,
    64'h00000000b06510eb,
    64'h00000000547aff27,
    64'h00000000bbaef3b2,
    64'h000000001608d275
};

localparam [63:0] WBL_ROM9 [0:63] = '{
    64'hff66789fbacd0963,
    64'hb33ccfa6780c837c,
    64'hd2e8df0025132c77,
    64'h000000002eec1a7b,
    64'h000000001c5f1bf2,
    64'h00000000a6976e6b,
    64'h00000000b4445a6f,
    64'h00000000c617a0c5,
    64'h00000000e8c45230,
    64'h00000000dda73b01,
    64'h00000000747ed667,
    64'h000000001f3db32b,
    64'h000000004b6429fe,
    64'h00000000bd5de3d7,
    64'h000000008b192fab,
    64'h000000008a738476,
    64'h00000000706053ca,
    64'h000000003e81d182,
    64'h00000000b54f00c9,
    64'h0000000066dced7d,
    64'h00000000482220fa,
    64'h00000000032afc59,
    64'h00000000f690b147,
    64'h000000000e885bf0,
    64'h0000000061466aad,
    64'h0000000035eecbd4,
    64'h0000000057b8bea2,
    64'h00000000b91439af,
    64'h0000000086de4a9c,
    64'h00000000c15e4ca4,
    64'h000000001d0b5872,
    64'h000000009edbcfc0,
    64'h00998760e1e0d0b7,
    64'h4cc33059f832effd,
    64'h2d172000983aaa93,
    64'h00000000110afb26,
    64'h0000000069494336,
    64'h00000000d9064d3f,
    64'h000000008e2433f7,
    64'h00000000945c85cc,
    64'h000000009bc24534,
    64'h000000001ed3f9a5,
    64'h0000000087ac02e5,
    64'h00000000e9627ff1,
    64'h00000000ce915071,
    64'h0000000055953cd8,
    64'h0000000028e49f31,
    64'h00000000df79a815,
    64'h000000008ce75104,
    64'h00000000a1c8a3c7,
    64'h0000000089374023,
    64'h000000000d6d8fc3,
    64'h00000000bf8d9218,
    64'h00000000e6d59d96,
    64'h00000000424e3805,
    64'h0000000068a9f59a,
    64'h00000000416cbc07,
    64'h000000009956b612,
    64'h000000002df4da80,
    64'h000000000fea21e2,
    64'h00000000b06510eb,
    64'h00000000547aff27,
    64'h00000000bbaef3b2,
    64'h000000001608d275
};

localparam [63:0] WBL_ROM10 [0:63] = '{
    64'h55bbc9f4bacd0963,
    64'h90bf3369780c837c,
    64'h8b095e0025132c77,
    64'h000000002eec1a7b,
    64'h000000001c5f1bf2,
    64'h00000000a6976e6b,
    64'h00000000b4445a6f,
    64'h00000000c617a0c5,
    64'h00000000e8c45230,
    64'h00000000dda73b01,
    64'h00000000747ed667,
    64'h000000001f3db32b,
    64'h000000004b6429fe,
    64'h00000000bd5de3d7,
    64'h000000008b192fab,
    64'h000000008a738476,
    64'h00000000706053ca,
    64'h000000003e81d182,
    64'h00000000b54f00c9,
    64'h0000000066dced7d,
    64'h00000000482220fa,
    64'h00000000032afc59,
    64'h00000000f690b147,
    64'h000000000e885bf0,
    64'h0000000061466aad,
    64'h0000000035eecbd4,
    64'h0000000057b8bea2,
    64'h00000000b91439af,
    64'h0000000086de4a9c,
    64'h00000000c15e4ca4,
    64'h000000001d0b5872,
    64'h000000009edbcfc0,
    64'haa44360be1e0d0b7,
    64'h6f40cc96f832effd,
    64'h74f6a100983aaa93,
    64'h00000000110afb26,
    64'h0000000069494336,
    64'h00000000d9064d3f,
    64'h000000008e2433f7,
    64'h00000000945c85cc,
    64'h000000009bc24534,
    64'h000000001ed3f9a5,
    64'h0000000087ac02e5,
    64'h00000000e9627ff1,
    64'h00000000ce915071,
    64'h0000000055953cd8,
    64'h0000000028e49f31,
    64'h00000000df79a815,
    64'h000000008ce75104,
    64'h00000000a1c8a3c7,
    64'h0000000089374023,
    64'h000000000d6d8fc3,
    64'h00000000bf8d9218,
    64'h00000000e6d59d96,
    64'h00000000424e3805,
    64'h0000000068a9f59a,
    64'h00000000416cbc07,
    64'h000000009956b612,
    64'h000000002df4da80,
    64'h000000000fea21e2,
    64'h00000000b06510eb,
    64'h00000000547aff27,
    64'h00000000bbaef3b2,
    64'h000000001608d275
};

localparam [63:0] WBL_ROM11 [0:63] = '{
    64'h336921d4bacd0963,
    64'hef267835780c837c,
    64'h6e27790025132c77,
    64'h000000002eec1a7b,
    64'h000000001c5f1bf2,
    64'h00000000a6976e6b,
    64'h00000000b4445a6f,
    64'h00000000c617a0c5,
    64'h00000000e8c45230,
    64'h00000000dda73b01,
    64'h00000000747ed667,
    64'h000000001f3db32b,
    64'h000000004b6429fe,
    64'h00000000bd5de3d7,
    64'h000000008b192fab,
    64'h000000008a738476,
    64'h00000000706053ca,
    64'h000000003e81d182,
    64'h00000000b54f00c9,
    64'h0000000066dced7d,
    64'h00000000482220fa,
    64'h00000000032afc59,
    64'h00000000f690b147,
    64'h000000000e885bf0,
    64'h0000000061466aad,
    64'h0000000035eecbd4,
    64'h0000000057b8bea2,
    64'h00000000b91439af,
    64'h0000000086de4a9c,
    64'h00000000c15e4ca4,
    64'h000000001d0b5872,
    64'h000000009edbcfc0,
    64'hcc96de2be1e0d0b7,
    64'h10d987caf832effd,
    64'h91d88600983aaa93,
    64'h00000000110afb26,
    64'h0000000069494336,
    64'h00000000d9064d3f,
    64'h000000008e2433f7,
    64'h00000000945c85cc,
    64'h000000009bc24534,
    64'h000000001ed3f9a5,
    64'h0000000087ac02e5,
    64'h00000000e9627ff1,
    64'h00000000ce915071,
    64'h0000000055953cd8,
    64'h0000000028e49f31,
    64'h00000000df79a815,
    64'h000000008ce75104,
    64'h00000000a1c8a3c7,
    64'h0000000089374023,
    64'h000000000d6d8fc3,
    64'h00000000bf8d9218,
    64'h00000000e6d59d96,
    64'h00000000424e3805,
    64'h0000000068a9f59a,
    64'h00000000416cbc07,
    64'h000000009956b612,
    64'h000000002df4da80,
    64'h000000000fea21e2,
    64'h00000000b06510eb,
    64'h00000000547aff27,
    64'h00000000bbaef3b2,
    64'h000000001608d275
};

localparam [63:0] WBL_ROM12 [0:63] = '{
    64'h0ff369debacd0963,
    64'h4df1c1fe780c837c,
    64'h3297460025132c77,
    64'h000000002eec1a7b,
    64'h000000001c5f1bf2,
    64'h00000000a6976e6b,
    64'h00000000b4445a6f,
    64'h00000000c617a0c5,
    64'h00000000e8c45230,
    64'h00000000dda73b01,
    64'h00000000747ed667,
    64'h000000001f3db32b,
    64'h000000004b6429fe,
    64'h00000000bd5de3d7,
    64'h000000008b192fab,
    64'h000000008a738476,
    64'h00000000706053ca,
    64'h000000003e81d182,
    64'h00000000b54f00c9,
    64'h0000000066dced7d,
    64'h00000000482220fa,
    64'h00000000032afc59,
    64'h00000000f690b147,
    64'h000000000e885bf0,
    64'h0000000061466aad,
    64'h0000000035eecbd4,
    64'h0000000057b8bea2,
    64'h00000000b91439af,
    64'h0000000086de4a9c,
    64'h00000000c15e4ca4,
    64'h000000001d0b5872,
    64'h000000009edbcfc0,
    64'hf00c9621e1e0d0b7,
    64'hb20e3e01f832effd,
    64'hcd68b900983aaa93,
    64'h00000000110afb26,
    64'h0000000069494336,
    64'h00000000d9064d3f,
    64'h000000008e2433f7,
    64'h00000000945c85cc,
    64'h000000009bc24534,
    64'h000000001ed3f9a5,
    64'h0000000087ac02e5,
    64'h00000000e9627ff1,
    64'h00000000ce915071,
    64'h0000000055953cd8,
    64'h0000000028e49f31,
    64'h00000000df79a815,
    64'h000000008ce75104,
    64'h00000000a1c8a3c7,
    64'h0000000089374023,
    64'h000000000d6d8fc3,
    64'h00000000bf8d9218,
    64'h00000000e6d59d96,
    64'h00000000424e3805,
    64'h0000000068a9f59a,
    64'h00000000416cbc07,
    64'h000000009956b612,
    64'h000000002df4da80,
    64'h000000000fea21e2,
    64'h00000000b06510eb,
    64'h00000000547aff27,
    64'h00000000bbaef3b2,
    64'h000000001608d275
};

localparam [63:0] WBL_ROM13 [0:63] = '{
    64'h0055bb9cbacd0963,
    64'he52ed8e0780c837c,
    64'h7fccf00025132c77,
    64'h000000002eec1a7b,
    64'h000000001c5f1bf2,
    64'h00000000a6976e6b,
    64'h00000000b4445a6f,
    64'h00000000c617a0c5,
    64'h00000000e8c45230,
    64'h00000000dda73b01,
    64'h00000000747ed667,
    64'h000000001f3db32b,
    64'h000000004b6429fe,
    64'h00000000bd5de3d7,
    64'h000000008b192fab,
    64'h000000008a738476,
    64'h00000000706053ca,
    64'h000000003e81d182,
    64'h00000000b54f00c9,
    64'h0000000066dced7d,
    64'h00000000482220fa,
    64'h00000000032afc59,
    64'h00000000f690b147,
    64'h000000000e885bf0,
    64'h0000000061466aad,
    64'h0000000035eecbd4,
    64'h0000000057b8bea2,
    64'h00000000b91439af,
    64'h0000000086de4a9c,
    64'h00000000c15e4ca4,
    64'h000000001d0b5872,
    64'h000000009edbcfc0,
    64'hffaa4463e1e0d0b7,
    64'h1ad1271ff832effd,
    64'h80330f00983aaa93,
    64'h00000000110afb26,
    64'h0000000069494336,
    64'h00000000d9064d3f,
    64'h000000008e2433f7,
    64'h00000000945c85cc,
    64'h000000009bc24534,
    64'h000000001ed3f9a5,
    64'h0000000087ac02e5,
    64'h00000000e9627ff1,
    64'h00000000ce915071,
    64'h0000000055953cd8,
    64'h0000000028e49f31,
    64'h00000000df79a815,
    64'h000000008ce75104,
    64'h00000000a1c8a3c7,
    64'h0000000089374023,
    64'h000000000d6d8fc3,
    64'h00000000bf8d9218,
    64'h00000000e6d59d96,
    64'h00000000424e3805,
    64'h0000000068a9f59a,
    64'h00000000416cbc07,
    64'h000000009956b612,
    64'h000000002df4da80,
    64'h000000000fea21e2,
    64'h00000000b06510eb,
    64'h00000000547aff27,
    64'h00000000bbaef3b2,
    64'h000000001608d275
};

localparam [63:0] WBL_ROM14 [0:63] = '{
    64'h00ff3396bacd0963,
    64'heddbe383780c837c,
    64'h5612420025132c77,
    64'h000000002eec1a7b,
    64'h000000001c5f1bf2,
    64'h00000000a6976e6b,
    64'h00000000b4445a6f,
    64'h00000000c617a0c5,
    64'h00000000e8c45230,
    64'h00000000dda73b01,
    64'h00000000747ed667,
    64'h000000001f3db32b,
    64'h000000004b6429fe,
    64'h00000000bd5de3d7,
    64'h000000008b192fab,
    64'h000000008a738476,
    64'h00000000706053ca,
    64'h000000003e81d182,
    64'h00000000b54f00c9,
    64'h0000000066dced7d,
    64'h00000000482220fa,
    64'h00000000032afc59,
    64'h00000000f690b147,
    64'h000000000e885bf0,
    64'h0000000061466aad,
    64'h0000000035eecbd4,
    64'h0000000057b8bea2,
    64'h00000000b91439af,
    64'h0000000086de4a9c,
    64'h00000000c15e4ca4,
    64'h000000001d0b5872,
    64'h000000009edbcfc0,
    64'hff00cc69e1e0d0b7,
    64'h12241c7cf832effd,
    64'ha9edbd00983aaa93,
    64'h00000000110afb26,
    64'h0000000069494336,
    64'h00000000d9064d3f,
    64'h000000008e2433f7,
    64'h00000000945c85cc,
    64'h000000009bc24534,
    64'h000000001ed3f9a5,
    64'h0000000087ac02e5,
    64'h00000000e9627ff1,
    64'h00000000ce915071,
    64'h0000000055953cd8,
    64'h0000000028e49f31,
    64'h00000000df79a815,
    64'h000000008ce75104,
    64'h00000000a1c8a3c7,
    64'h0000000089374023,
    64'h000000000d6d8fc3,
    64'h00000000bf8d9218,
    64'h00000000e6d59d96,
    64'h00000000424e3805,
    64'h0000000068a9f59a,
    64'h00000000416cbc07,
    64'h000000009956b612,
    64'h000000002df4da80,
    64'h000000000fea21e2,
    64'h00000000b06510eb,
    64'h00000000547aff27,
    64'h00000000bbaef3b2,
    64'h000000001608d275
};

localparam [63:0] WBL_ROM15 [0:63] = '{
    64'h005511ebbacd0963,
    64'h895e4da4780c837c,
    64'h8551410025132c77,
    64'h000000002eec1a7b,
    64'h000000001c5f1bf2,
    64'h00000000a6976e6b,
    64'h00000000b4445a6f,
    64'h00000000c617a0c5,
    64'h00000000e8c45230,
    64'h00000000dda73b01,
    64'h00000000747ed667,
    64'h000000001f3db32b,
    64'h000000004b6429fe,
    64'h00000000bd5de3d7,
    64'h000000008b192fab,
    64'h000000008a738476,
    64'h00000000706053ca,
    64'h000000003e81d182,
    64'h00000000b54f00c9,
    64'h0000000066dced7d,
    64'h00000000482220fa,
    64'h00000000032afc59,
    64'h00000000f690b147,
    64'h000000000e885bf0,
    64'h0000000061466aad,
    64'h0000000035eecbd4,
    64'h0000000057b8bea2,
    64'h00000000b91439af,
    64'h0000000086de4a9c,
    64'h00000000c15e4ca4,
    64'h000000001d0b5872,
    64'h000000009edbcfc0,
    64'hffaaee14e1e0d0b7,
    64'h76a1b25bf832effd,
    64'h7aaebe00983aaa93,
    64'h00000000110afb26,
    64'h0000000069494336,
    64'h00000000d9064d3f,
    64'h000000008e2433f7,
    64'h00000000945c85cc,
    64'h000000009bc24534,
    64'h000000001ed3f9a5,
    64'h0000000087ac02e5,
    64'h00000000e9627ff1,
    64'h00000000ce915071,
    64'h0000000055953cd8,
    64'h0000000028e49f31,
    64'h00000000df79a815,
    64'h000000008ce75104,
    64'h00000000a1c8a3c7,
    64'h0000000089374023,
    64'h000000000d6d8fc3,
    64'h00000000bf8d9218,
    64'h00000000e6d59d96,
    64'h00000000424e3805,
    64'h0000000068a9f59a,
    64'h00000000416cbc07,
    64'h000000009956b612,
    64'h000000002df4da80,
    64'h000000000fea21e2,
    64'h00000000b06510eb,
    64'h00000000547aff27,
    64'h00000000bbaef3b2,
    64'h000000001608d275
};

localparam [63:0] WBL_ROM16 [0:63] = '{
    64'h00ff99b4bacd0963,
    64'hc5fb3692780c837c,
    64'h17ec250025132c77,
    64'h000000002eec1a7b,
    64'h000000001c5f1bf2,
    64'h00000000a6976e6b,
    64'h00000000b4445a6f,
    64'h00000000c617a0c5,
    64'h00000000e8c45230,
    64'h00000000dda73b01,
    64'h00000000747ed667,
    64'h000000001f3db32b,
    64'h000000004b6429fe,
    64'h00000000bd5de3d7,
    64'h000000008b192fab,
    64'h000000008a738476,
    64'h00000000706053ca,
    64'h000000003e81d182,
    64'h00000000b54f00c9,
    64'h0000000066dced7d,
    64'h00000000482220fa,
    64'h00000000032afc59,
    64'h00000000f690b147,
    64'h000000000e885bf0,
    64'h0000000061466aad,
    64'h0000000035eecbd4,
    64'h0000000057b8bea2,
    64'h00000000b91439af,
    64'h0000000086de4a9c,
    64'h00000000c15e4ca4,
    64'h000000001d0b5872,
    64'h000000009edbcfc0,
    64'hff00664be1e0d0b7,
    64'h3a04c96df832effd,
    64'he813da00983aaa93,
    64'h00000000110afb26,
    64'h0000000069494336,
    64'h00000000d9064d3f,
    64'h000000008e2433f7,
    64'h00000000945c85cc,
    64'h000000009bc24534,
    64'h000000001ed3f9a5,
    64'h0000000087ac02e5,
    64'h00000000e9627ff1,
    64'h00000000ce915071,
    64'h0000000055953cd8,
    64'h0000000028e49f31,
    64'h00000000df79a815,
    64'h000000008ce75104,
    64'h00000000a1c8a3c7,
    64'h0000000089374023,
    64'h000000000d6d8fc3,
    64'h00000000bf8d9218,
    64'h00000000e6d59d96,
    64'h00000000424e3805,
    64'h0000000068a9f59a,
    64'h00000000416cbc07,
    64'h000000009956b612,
    64'h000000002df4da80,
    64'h000000000fea21e2,
    64'h00000000b06510eb,
    64'h00000000547aff27,
    64'h00000000bbaef3b2,
    64'h000000001608d275
};

