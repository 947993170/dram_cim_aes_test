wire [63:0] WBL_ROM1 [0:63];
assign WBL_ROM1[0] = 64'h00005511bacd0963;
assign WBL_ROM1[1] = 64'heb766d24780c837c;
assign WBL_ROM1[2] = 64'hd015ee0025132c77;
assign WBL_ROM1[3] = 64'h000000002eec1a7b;
assign WBL_ROM1[4] = 64'h000000001c5f1bf2;
assign WBL_ROM1[5] = 64'h00000000a6976e6b;
assign WBL_ROM1[6] = 64'h00000000b4445a6f;
assign WBL_ROM1[7] = 64'h00000000c617a0c5;
assign WBL_ROM1[8] = 64'h00000000e8c45230;
assign WBL_ROM1[9] = 64'h00000000dda73b01;
assign WBL_ROM1[10] = 64'h00000000747ed667;
assign WBL_ROM1[11] = 64'h000000001f3db32b;
assign WBL_ROM1[12] = 64'h000000004b6429fe;
assign WBL_ROM1[13] = 64'h00000000bd5de3d7;
assign WBL_ROM1[14] = 64'h000000008b192fab;
assign WBL_ROM1[15] = 64'h000000008a738476;
assign WBL_ROM1[16] = 64'h00000000706053ca;
assign WBL_ROM1[17] = 64'h000000003e81d182;
assign WBL_ROM1[18] = 64'h00000000b54f00c9;
assign WBL_ROM1[19] = 64'h0000000066dced7d;
assign WBL_ROM1[20] = 64'h00000000482220fa;
assign WBL_ROM1[21] = 64'h00000000032afc59;
assign WBL_ROM1[22] = 64'h00000000f690b147;
assign WBL_ROM1[23] = 64'h000000000e885bf0;
assign WBL_ROM1[24] = 64'h0000000061466aad;
assign WBL_ROM1[25] = 64'h0000000035eecbd4;
assign WBL_ROM1[26] = 64'h0000000057b8bea2;
assign WBL_ROM1[27] = 64'h00000000b91439af;
assign WBL_ROM1[28] = 64'h0000000086de4a9c;
assign WBL_ROM1[29] = 64'h00000000c15e4ca4;
assign WBL_ROM1[30] = 64'h000000001d0b5872;
assign WBL_ROM1[31] = 64'h000000009edbcfc0;
assign WBL_ROM1[32] = 64'hffffaaeee1e0d0b7;
assign WBL_ROM1[33] = 64'h148992dbf832effd;
assign WBL_ROM1[34] = 64'h2fea1100983aaa93;
assign WBL_ROM1[35] = 64'h00000000110afb26;
assign WBL_ROM1[36] = 64'h0000000069494336;
assign WBL_ROM1[37] = 64'h00000000d9064d3f;
assign WBL_ROM1[38] = 64'h000000008e2433f7;
assign WBL_ROM1[39] = 64'h00000000945c85cc;
assign WBL_ROM1[40] = 64'h000000009bc24534;
assign WBL_ROM1[41] = 64'h000000001ed3f9a5;
assign WBL_ROM1[42] = 64'h0000000087ac02e5;
assign WBL_ROM1[43] = 64'h00000000e9627ff1;
assign WBL_ROM1[44] = 64'h00000000ce915071;
assign WBL_ROM1[45] = 64'h0000000055953cd8;
assign WBL_ROM1[46] = 64'h0000000028e49f31;
assign WBL_ROM1[47] = 64'h00000000df79a815;
assign WBL_ROM1[48] = 64'h000000008ce75104;
assign WBL_ROM1[49] = 64'h00000000a1c8a3c7;
assign WBL_ROM1[50] = 64'h0000000089374023;
assign WBL_ROM1[51] = 64'h000000000d6d8fc3;
assign WBL_ROM1[52] = 64'h00000000bf8d9218;
assign WBL_ROM1[53] = 64'h00000000e6d59d96;
assign WBL_ROM1[54] = 64'h00000000424e3805;
assign WBL_ROM1[55] = 64'h0000000068a9f59a;
assign WBL_ROM1[56] = 64'h00000000416cbc07;
assign WBL_ROM1[57] = 64'h000000009956b612;
assign WBL_ROM1[58] = 64'h000000002df4da80;
assign WBL_ROM1[59] = 64'h000000000fea21e2;
assign WBL_ROM1[60] = 64'h00000000b06510eb;
assign WBL_ROM1[61] = 64'h00000000547aff27;
assign WBL_ROM1[62] = 64'h00000000bbaef3b2;
assign WBL_ROM1[63] = 64'h000000001608d275;

wire [63:0] WBL_ROM2 [0:63];
assign WBL_ROM2[0] = 64'h55bbc9a1bacd0963;
assign WBL_ROM2[1] = 64'hd445fb36780c837c;
assign WBL_ROM2[2] = 64'hc753bc0025132c77;
assign WBL_ROM2[3] = 64'h000000002eec1a7b;
assign WBL_ROM2[4] = 64'h000000001c5f1bf2;
assign WBL_ROM2[5] = 64'h00000000a6976e6b;
assign WBL_ROM2[6] = 64'h00000000b4445a6f;
assign WBL_ROM2[7] = 64'h00000000c617a0c5;
assign WBL_ROM2[8] = 64'h00000000e8c45230;
assign WBL_ROM2[9] = 64'h00000000dda73b01;
assign WBL_ROM2[10] = 64'h00000000747ed667;
assign WBL_ROM2[11] = 64'h000000001f3db32b;
assign WBL_ROM2[12] = 64'h000000004b6429fe;
assign WBL_ROM2[13] = 64'h00000000bd5de3d7;
assign WBL_ROM2[14] = 64'h000000008b192fab;
assign WBL_ROM2[15] = 64'h000000008a738476;
assign WBL_ROM2[16] = 64'h00000000706053ca;
assign WBL_ROM2[17] = 64'h000000003e81d182;
assign WBL_ROM2[18] = 64'h00000000b54f00c9;
assign WBL_ROM2[19] = 64'h0000000066dced7d;
assign WBL_ROM2[20] = 64'h00000000482220fa;
assign WBL_ROM2[21] = 64'h00000000032afc59;
assign WBL_ROM2[22] = 64'h00000000f690b147;
assign WBL_ROM2[23] = 64'h000000000e885bf0;
assign WBL_ROM2[24] = 64'h0000000061466aad;
assign WBL_ROM2[25] = 64'h0000000035eecbd4;
assign WBL_ROM2[26] = 64'h0000000057b8bea2;
assign WBL_ROM2[27] = 64'h00000000b91439af;
assign WBL_ROM2[28] = 64'h0000000086de4a9c;
assign WBL_ROM2[29] = 64'h00000000c15e4ca4;
assign WBL_ROM2[30] = 64'h000000001d0b5872;
assign WBL_ROM2[31] = 64'h000000009edbcfc0;
assign WBL_ROM2[32] = 64'haa44365ee1e0d0b7;
assign WBL_ROM2[33] = 64'h2bba04c9f832effd;
assign WBL_ROM2[34] = 64'h38ac4300983aaa93;
assign WBL_ROM2[35] = 64'h00000000110afb26;
assign WBL_ROM2[36] = 64'h0000000069494336;
assign WBL_ROM2[37] = 64'h00000000d9064d3f;
assign WBL_ROM2[38] = 64'h000000008e2433f7;
assign WBL_ROM2[39] = 64'h00000000945c85cc;
assign WBL_ROM2[40] = 64'h000000009bc24534;
assign WBL_ROM2[41] = 64'h000000001ed3f9a5;
assign WBL_ROM2[42] = 64'h0000000087ac02e5;
assign WBL_ROM2[43] = 64'h00000000e9627ff1;
assign WBL_ROM2[44] = 64'h00000000ce915071;
assign WBL_ROM2[45] = 64'h0000000055953cd8;
assign WBL_ROM2[46] = 64'h0000000028e49f31;
assign WBL_ROM2[47] = 64'h00000000df79a815;
assign WBL_ROM2[48] = 64'h000000008ce75104;
assign WBL_ROM2[49] = 64'h00000000a1c8a3c7;
assign WBL_ROM2[50] = 64'h0000000089374023;
assign WBL_ROM2[51] = 64'h000000000d6d8fc3;
assign WBL_ROM2[52] = 64'h00000000bf8d9218;
assign WBL_ROM2[53] = 64'h00000000e6d59d96;
assign WBL_ROM2[54] = 64'h00000000424e3805;
assign WBL_ROM2[55] = 64'h0000000068a9f59a;
assign WBL_ROM2[56] = 64'h00000000416cbc07;
assign WBL_ROM2[57] = 64'h000000009956b612;
assign WBL_ROM2[58] = 64'h000000002df4da80;
assign WBL_ROM2[59] = 64'h000000000fea21e2;
assign WBL_ROM2[60] = 64'h00000000b06510eb;
assign WBL_ROM2[61] = 64'h00000000547aff27;
assign WBL_ROM2[62] = 64'h00000000bbaef3b2;
assign WBL_ROM2[63] = 64'h000000001608d275;

wire [63:0] WBL_ROM3 [0:63];
assign WBL_ROM3[0] = 64'h33c3fccfbacd0963;
assign WBL_ROM3[1] = 64'hf396ed8e780c837c;
assign WBL_ROM3[2] = 64'hf297460025132c77;
assign WBL_ROM3[3] = 64'h000000002eec1a7b;
assign WBL_ROM3[4] = 64'h000000001c5f1bf2;
assign WBL_ROM3[5] = 64'h00000000a6976e6b;
assign WBL_ROM3[6] = 64'h00000000b4445a6f;
assign WBL_ROM3[7] = 64'h00000000c617a0c5;
assign WBL_ROM3[8] = 64'h00000000e8c45230;
assign WBL_ROM3[9] = 64'h00000000dda73b01;
assign WBL_ROM3[10] = 64'h00000000747ed667;
assign WBL_ROM3[11] = 64'h000000001f3db32b;
assign WBL_ROM3[12] = 64'h000000004b6429fe;
assign WBL_ROM3[13] = 64'h00000000bd5de3d7;
assign WBL_ROM3[14] = 64'h000000008b192fab;
assign WBL_ROM3[15] = 64'h000000008a738476;
assign WBL_ROM3[16] = 64'h00000000706053ca;
assign WBL_ROM3[17] = 64'h000000003e81d182;
assign WBL_ROM3[18] = 64'h00000000b54f00c9;
assign WBL_ROM3[19] = 64'h0000000066dced7d;
assign WBL_ROM3[20] = 64'h00000000482220fa;
assign WBL_ROM3[21] = 64'h00000000032afc59;
assign WBL_ROM3[22] = 64'h00000000f690b147;
assign WBL_ROM3[23] = 64'h000000000e885bf0;
assign WBL_ROM3[24] = 64'h0000000061466aad;
assign WBL_ROM3[25] = 64'h0000000035eecbd4;
assign WBL_ROM3[26] = 64'h0000000057b8bea2;
assign WBL_ROM3[27] = 64'h00000000b91439af;
assign WBL_ROM3[28] = 64'h0000000086de4a9c;
assign WBL_ROM3[29] = 64'h00000000c15e4ca4;
assign WBL_ROM3[30] = 64'h000000001d0b5872;
assign WBL_ROM3[31] = 64'h000000009edbcfc0;
assign WBL_ROM3[32] = 64'hcc3c0330e1e0d0b7;
assign WBL_ROM3[33] = 64'h0c691271f832effd;
assign WBL_ROM3[34] = 64'h0d68b900983aaa93;
assign WBL_ROM3[35] = 64'h00000000110afb26;
assign WBL_ROM3[36] = 64'h0000000069494336;
assign WBL_ROM3[37] = 64'h00000000d9064d3f;
assign WBL_ROM3[38] = 64'h000000008e2433f7;
assign WBL_ROM3[39] = 64'h00000000945c85cc;
assign WBL_ROM3[40] = 64'h000000009bc24534;
assign WBL_ROM3[41] = 64'h000000001ed3f9a5;
assign WBL_ROM3[42] = 64'h0000000087ac02e5;
assign WBL_ROM3[43] = 64'h00000000e9627ff1;
assign WBL_ROM3[44] = 64'h00000000ce915071;
assign WBL_ROM3[45] = 64'h0000000055953cd8;
assign WBL_ROM3[46] = 64'h0000000028e49f31;
assign WBL_ROM3[47] = 64'h00000000df79a815;
assign WBL_ROM3[48] = 64'h000000008ce75104;
assign WBL_ROM3[49] = 64'h00000000a1c8a3c7;
assign WBL_ROM3[50] = 64'h0000000089374023;
assign WBL_ROM3[51] = 64'h000000000d6d8fc3;
assign WBL_ROM3[52] = 64'h00000000bf8d9218;
assign WBL_ROM3[53] = 64'h00000000e6d59d96;
assign WBL_ROM3[54] = 64'h00000000424e3805;
assign WBL_ROM3[55] = 64'h0000000068a9f59a;
assign WBL_ROM3[56] = 64'h00000000416cbc07;
assign WBL_ROM3[57] = 64'h000000009956b612;
assign WBL_ROM3[58] = 64'h000000002df4da80;
assign WBL_ROM3[59] = 64'h000000000fea21e2;
assign WBL_ROM3[60] = 64'h00000000b06510eb;
assign WBL_ROM3[61] = 64'h00000000547aff27;
assign WBL_ROM3[62] = 64'h00000000bbaef3b2;
assign WBL_ROM3[63] = 64'h000000001608d275;

wire [63:0] WBL_ROM4 [0:63];
assign WBL_ROM4[0] = 64'h0f0c5a1dbacd0963;
assign WBL_ROM4[1] = 64'h1bb6c706780c837c;
assign WBL_ROM4[2] = 64'h0706520025132c77;
assign WBL_ROM4[3] = 64'h000000002eec1a7b;
assign WBL_ROM4[4] = 64'h000000001c5f1bf2;
assign WBL_ROM4[5] = 64'h00000000a6976e6b;
assign WBL_ROM4[6] = 64'h00000000b4445a6f;
assign WBL_ROM4[7] = 64'h00000000c617a0c5;
assign WBL_ROM4[8] = 64'h00000000e8c45230;
assign WBL_ROM4[9] = 64'h00000000dda73b01;
assign WBL_ROM4[10] = 64'h00000000747ed667;
assign WBL_ROM4[11] = 64'h000000001f3db32b;
assign WBL_ROM4[12] = 64'h000000004b6429fe;
assign WBL_ROM4[13] = 64'h00000000bd5de3d7;
assign WBL_ROM4[14] = 64'h000000008b192fab;
assign WBL_ROM4[15] = 64'h000000008a738476;
assign WBL_ROM4[16] = 64'h00000000706053ca;
assign WBL_ROM4[17] = 64'h000000003e81d182;
assign WBL_ROM4[18] = 64'h00000000b54f00c9;
assign WBL_ROM4[19] = 64'h0000000066dced7d;
assign WBL_ROM4[20] = 64'h00000000482220fa;
assign WBL_ROM4[21] = 64'h00000000032afc59;
assign WBL_ROM4[22] = 64'h00000000f690b147;
assign WBL_ROM4[23] = 64'h000000000e885bf0;
assign WBL_ROM4[24] = 64'h0000000061466aad;
assign WBL_ROM4[25] = 64'h0000000035eecbd4;
assign WBL_ROM4[26] = 64'h0000000057b8bea2;
assign WBL_ROM4[27] = 64'h00000000b91439af;
assign WBL_ROM4[28] = 64'h0000000086de4a9c;
assign WBL_ROM4[29] = 64'h00000000c15e4ca4;
assign WBL_ROM4[30] = 64'h000000001d0b5872;
assign WBL_ROM4[31] = 64'h000000009edbcfc0;
assign WBL_ROM4[32] = 64'hf0f3a5e2e1e0d0b7;
assign WBL_ROM4[33] = 64'he44938f9f832effd;
assign WBL_ROM4[34] = 64'hf8f9ad00983aaa93;
assign WBL_ROM4[35] = 64'h00000000110afb26;
assign WBL_ROM4[36] = 64'h0000000069494336;
assign WBL_ROM4[37] = 64'h00000000d9064d3f;
assign WBL_ROM4[38] = 64'h000000008e2433f7;
assign WBL_ROM4[39] = 64'h00000000945c85cc;
assign WBL_ROM4[40] = 64'h000000009bc24534;
assign WBL_ROM4[41] = 64'h000000001ed3f9a5;
assign WBL_ROM4[42] = 64'h0000000087ac02e5;
assign WBL_ROM4[43] = 64'h00000000e9627ff1;
assign WBL_ROM4[44] = 64'h00000000ce915071;
assign WBL_ROM4[45] = 64'h0000000055953cd8;
assign WBL_ROM4[46] = 64'h0000000028e49f31;
assign WBL_ROM4[47] = 64'h00000000df79a815;
assign WBL_ROM4[48] = 64'h000000008ce75104;
assign WBL_ROM4[49] = 64'h00000000a1c8a3c7;
assign WBL_ROM4[50] = 64'h0000000089374023;
assign WBL_ROM4[51] = 64'h000000000d6d8fc3;
assign WBL_ROM4[52] = 64'h00000000bf8d9218;
assign WBL_ROM4[53] = 64'h00000000e6d59d96;
assign WBL_ROM4[54] = 64'h00000000424e3805;
assign WBL_ROM4[55] = 64'h0000000068a9f59a;
assign WBL_ROM4[56] = 64'h00000000416cbc07;
assign WBL_ROM4[57] = 64'h000000009956b612;
assign WBL_ROM4[58] = 64'h000000002df4da80;
assign WBL_ROM4[59] = 64'h000000000fea21e2;
assign WBL_ROM4[60] = 64'h00000000b06510eb;
assign WBL_ROM4[61] = 64'h00000000547aff27;
assign WBL_ROM4[62] = 64'h00000000bbaef3b2;
assign WBL_ROM4[63] = 64'h000000001608d275;

wire [63:0] WBL_ROM5 [0:63];
assign WBL_ROM5[0] = 64'h00ff99e1bacd0963;
assign WBL_ROM5[1] = 64'h7e98b5c4780c837c;
assign WBL_ROM5[2] = 64'h05fbc90025132c77;
assign WBL_ROM5[3] = 64'h000000002eec1a7b;
assign WBL_ROM5[4] = 64'h000000001c5f1bf2;
assign WBL_ROM5[5] = 64'h00000000a6976e6b;
assign WBL_ROM5[6] = 64'h00000000b4445a6f;
assign WBL_ROM5[7] = 64'h00000000c617a0c5;
assign WBL_ROM5[8] = 64'h00000000e8c45230;
assign WBL_ROM5[9] = 64'h00000000dda73b01;
assign WBL_ROM5[10] = 64'h00000000747ed667;
assign WBL_ROM5[11] = 64'h000000001f3db32b;
assign WBL_ROM5[12] = 64'h000000004b6429fe;
assign WBL_ROM5[13] = 64'h00000000bd5de3d7;
assign WBL_ROM5[14] = 64'h000000008b192fab;
assign WBL_ROM5[15] = 64'h000000008a738476;
assign WBL_ROM5[16] = 64'h00000000706053ca;
assign WBL_ROM5[17] = 64'h000000003e81d182;
assign WBL_ROM5[18] = 64'h00000000b54f00c9;
assign WBL_ROM5[19] = 64'h0000000066dced7d;
assign WBL_ROM5[20] = 64'h00000000482220fa;
assign WBL_ROM5[21] = 64'h00000000032afc59;
assign WBL_ROM5[22] = 64'h00000000f690b147;
assign WBL_ROM5[23] = 64'h000000000e885bf0;
assign WBL_ROM5[24] = 64'h0000000061466aad;
assign WBL_ROM5[25] = 64'h0000000035eecbd4;
assign WBL_ROM5[26] = 64'h0000000057b8bea2;
assign WBL_ROM5[27] = 64'h00000000b91439af;
assign WBL_ROM5[28] = 64'h0000000086de4a9c;
assign WBL_ROM5[29] = 64'h00000000c15e4ca4;
assign WBL_ROM5[30] = 64'h000000001d0b5872;
assign WBL_ROM5[31] = 64'h000000009edbcfc0;
assign WBL_ROM5[32] = 64'hff00661ee1e0d0b7;
assign WBL_ROM5[33] = 64'h81674a3bf832effd;
assign WBL_ROM5[34] = 64'hfa043600983aaa93;
assign WBL_ROM5[35] = 64'h00000000110afb26;
assign WBL_ROM5[36] = 64'h0000000069494336;
assign WBL_ROM5[37] = 64'h00000000d9064d3f;
assign WBL_ROM5[38] = 64'h000000008e2433f7;
assign WBL_ROM5[39] = 64'h00000000945c85cc;
assign WBL_ROM5[40] = 64'h000000009bc24534;
assign WBL_ROM5[41] = 64'h000000001ed3f9a5;
assign WBL_ROM5[42] = 64'h0000000087ac02e5;
assign WBL_ROM5[43] = 64'h00000000e9627ff1;
assign WBL_ROM5[44] = 64'h00000000ce915071;
assign WBL_ROM5[45] = 64'h0000000055953cd8;
assign WBL_ROM5[46] = 64'h0000000028e49f31;
assign WBL_ROM5[47] = 64'h00000000df79a815;
assign WBL_ROM5[48] = 64'h000000008ce75104;
assign WBL_ROM5[49] = 64'h00000000a1c8a3c7;
assign WBL_ROM5[50] = 64'h0000000089374023;
assign WBL_ROM5[51] = 64'h000000000d6d8fc3;
assign WBL_ROM5[52] = 64'h00000000bf8d9218;
assign WBL_ROM5[53] = 64'h00000000e6d59d96;
assign WBL_ROM5[54] = 64'h00000000424e3805;
assign WBL_ROM5[55] = 64'h0000000068a9f59a;
assign WBL_ROM5[56] = 64'h00000000416cbc07;
assign WBL_ROM5[57] = 64'h000000009956b612;
assign WBL_ROM5[58] = 64'h000000002df4da80;
assign WBL_ROM5[59] = 64'h000000000fea21e2;
assign WBL_ROM5[60] = 64'h00000000b06510eb;
assign WBL_ROM5[61] = 64'h00000000547aff27;
assign WBL_ROM5[62] = 64'h00000000bbaef3b2;
assign WBL_ROM5[63] = 64'h000000001608d275;

wire [63:0] WBL_ROM6 [0:63];
assign WBL_ROM6[0] = 64'h0055bbc9bacd0963;
assign WBL_ROM6[1] = 64'h5ee72c70780c837c;
assign WBL_ROM6[2] = 64'h3f662d0025132c77;
assign WBL_ROM6[3] = 64'h000000002eec1a7b;
assign WBL_ROM6[4] = 64'h000000001c5f1bf2;
assign WBL_ROM6[5] = 64'h00000000a6976e6b;
assign WBL_ROM6[6] = 64'h00000000b4445a6f;
assign WBL_ROM6[7] = 64'h00000000c617a0c5;
assign WBL_ROM6[8] = 64'h00000000e8c45230;
assign WBL_ROM6[9] = 64'h00000000dda73b01;
assign WBL_ROM6[10] = 64'h00000000747ed667;
assign WBL_ROM6[11] = 64'h000000001f3db32b;
assign WBL_ROM6[12] = 64'h000000004b6429fe;
assign WBL_ROM6[13] = 64'h00000000bd5de3d7;
assign WBL_ROM6[14] = 64'h000000008b192fab;
assign WBL_ROM6[15] = 64'h000000008a738476;
assign WBL_ROM6[16] = 64'h00000000706053ca;
assign WBL_ROM6[17] = 64'h000000003e81d182;
assign WBL_ROM6[18] = 64'h00000000b54f00c9;
assign WBL_ROM6[19] = 64'h0000000066dced7d;
assign WBL_ROM6[20] = 64'h00000000482220fa;
assign WBL_ROM6[21] = 64'h00000000032afc59;
assign WBL_ROM6[22] = 64'h00000000f690b147;
assign WBL_ROM6[23] = 64'h000000000e885bf0;
assign WBL_ROM6[24] = 64'h0000000061466aad;
assign WBL_ROM6[25] = 64'h0000000035eecbd4;
assign WBL_ROM6[26] = 64'h0000000057b8bea2;
assign WBL_ROM6[27] = 64'h00000000b91439af;
assign WBL_ROM6[28] = 64'h0000000086de4a9c;
assign WBL_ROM6[29] = 64'h00000000c15e4ca4;
assign WBL_ROM6[30] = 64'h000000001d0b5872;
assign WBL_ROM6[31] = 64'h000000009edbcfc0;
assign WBL_ROM6[32] = 64'hffaa4436e1e0d0b7;
assign WBL_ROM6[33] = 64'ha118d38ff832effd;
assign WBL_ROM6[34] = 64'hc099d200983aaa93;
assign WBL_ROM6[35] = 64'h00000000110afb26;
assign WBL_ROM6[36] = 64'h0000000069494336;
assign WBL_ROM6[37] = 64'h00000000d9064d3f;
assign WBL_ROM6[38] = 64'h000000008e2433f7;
assign WBL_ROM6[39] = 64'h00000000945c85cc;
assign WBL_ROM6[40] = 64'h000000009bc24534;
assign WBL_ROM6[41] = 64'h000000001ed3f9a5;
assign WBL_ROM6[42] = 64'h0000000087ac02e5;
assign WBL_ROM6[43] = 64'h00000000e9627ff1;
assign WBL_ROM6[44] = 64'h00000000ce915071;
assign WBL_ROM6[45] = 64'h0000000055953cd8;
assign WBL_ROM6[46] = 64'h0000000028e49f31;
assign WBL_ROM6[47] = 64'h00000000df79a815;
assign WBL_ROM6[48] = 64'h000000008ce75104;
assign WBL_ROM6[49] = 64'h00000000a1c8a3c7;
assign WBL_ROM6[50] = 64'h0000000089374023;
assign WBL_ROM6[51] = 64'h000000000d6d8fc3;
assign WBL_ROM6[52] = 64'h00000000bf8d9218;
assign WBL_ROM6[53] = 64'h00000000e6d59d96;
assign WBL_ROM6[54] = 64'h00000000424e3805;
assign WBL_ROM6[55] = 64'h0000000068a9f59a;
assign WBL_ROM6[56] = 64'h00000000416cbc07;
assign WBL_ROM6[57] = 64'h000000009956b612;
assign WBL_ROM6[58] = 64'h000000002df4da80;
assign WBL_ROM6[59] = 64'h000000000fea21e2;
assign WBL_ROM6[60] = 64'h00000000b06510eb;
assign WBL_ROM6[61] = 64'h00000000547aff27;
assign WBL_ROM6[62] = 64'h00000000bbaef3b2;
assign WBL_ROM6[63] = 64'h000000001608d275;

wire [63:0] WBL_ROM7 [0:63];
assign WBL_ROM7[0] = 64'h00ff6678bacd0963;
assign WBL_ROM7[1] = 64'hca08a07f780c837c;
assign WBL_ROM7[2] = 64'h99b43a0025132c77;
assign WBL_ROM7[3] = 64'h000000002eec1a7b;
assign WBL_ROM7[4] = 64'h000000001c5f1bf2;
assign WBL_ROM7[5] = 64'h00000000a6976e6b;
assign WBL_ROM7[6] = 64'h00000000b4445a6f;
assign WBL_ROM7[7] = 64'h00000000c617a0c5;
assign WBL_ROM7[8] = 64'h00000000e8c45230;
assign WBL_ROM7[9] = 64'h00000000dda73b01;
assign WBL_ROM7[10] = 64'h00000000747ed667;
assign WBL_ROM7[11] = 64'h000000001f3db32b;
assign WBL_ROM7[12] = 64'h000000004b6429fe;
assign WBL_ROM7[13] = 64'h00000000bd5de3d7;
assign WBL_ROM7[14] = 64'h000000008b192fab;
assign WBL_ROM7[15] = 64'h000000008a738476;
assign WBL_ROM7[16] = 64'h00000000706053ca;
assign WBL_ROM7[17] = 64'h000000003e81d182;
assign WBL_ROM7[18] = 64'h00000000b54f00c9;
assign WBL_ROM7[19] = 64'h0000000066dced7d;
assign WBL_ROM7[20] = 64'h00000000482220fa;
assign WBL_ROM7[21] = 64'h00000000032afc59;
assign WBL_ROM7[22] = 64'h00000000f690b147;
assign WBL_ROM7[23] = 64'h000000000e885bf0;
assign WBL_ROM7[24] = 64'h0000000061466aad;
assign WBL_ROM7[25] = 64'h0000000035eecbd4;
assign WBL_ROM7[26] = 64'h0000000057b8bea2;
assign WBL_ROM7[27] = 64'h00000000b91439af;
assign WBL_ROM7[28] = 64'h0000000086de4a9c;
assign WBL_ROM7[29] = 64'h00000000c15e4ca4;
assign WBL_ROM7[30] = 64'h000000001d0b5872;
assign WBL_ROM7[31] = 64'h000000009edbcfc0;
assign WBL_ROM7[32] = 64'hff009987e1e0d0b7;
assign WBL_ROM7[33] = 64'h35f75f80f832effd;
assign WBL_ROM7[34] = 64'h664bc500983aaa93;
assign WBL_ROM7[35] = 64'h00000000110afb26;
assign WBL_ROM7[36] = 64'h0000000069494336;
assign WBL_ROM7[37] = 64'h00000000d9064d3f;
assign WBL_ROM7[38] = 64'h000000008e2433f7;
assign WBL_ROM7[39] = 64'h00000000945c85cc;
assign WBL_ROM7[40] = 64'h000000009bc24534;
assign WBL_ROM7[41] = 64'h000000001ed3f9a5;
assign WBL_ROM7[42] = 64'h0000000087ac02e5;
assign WBL_ROM7[43] = 64'h00000000e9627ff1;
assign WBL_ROM7[44] = 64'h00000000ce915071;
assign WBL_ROM7[45] = 64'h0000000055953cd8;
assign WBL_ROM7[46] = 64'h0000000028e49f31;
assign WBL_ROM7[47] = 64'h00000000df79a815;
assign WBL_ROM7[48] = 64'h000000008ce75104;
assign WBL_ROM7[49] = 64'h00000000a1c8a3c7;
assign WBL_ROM7[50] = 64'h0000000089374023;
assign WBL_ROM7[51] = 64'h000000000d6d8fc3;
assign WBL_ROM7[52] = 64'h00000000bf8d9218;
assign WBL_ROM7[53] = 64'h00000000e6d59d96;
assign WBL_ROM7[54] = 64'h00000000424e3805;
assign WBL_ROM7[55] = 64'h0000000068a9f59a;
assign WBL_ROM7[56] = 64'h00000000416cbc07;
assign WBL_ROM7[57] = 64'h000000009956b612;
assign WBL_ROM7[58] = 64'h000000002df4da80;
assign WBL_ROM7[59] = 64'h000000000fea21e2;
assign WBL_ROM7[60] = 64'h00000000b06510eb;
assign WBL_ROM7[61] = 64'h00000000547aff27;
assign WBL_ROM7[62] = 64'h00000000bbaef3b2;
assign WBL_ROM7[63] = 64'h000000001608d275;

wire [63:0] WBL_ROM8 [0:63];
assign WBL_ROM8[0] = 64'h00aaddb1bacd0963;
assign WBL_ROM8[1] = 64'h6b763835780c837c;
assign WBL_ROM8[2] = 64'h6e272c0025132c77;
assign WBL_ROM8[3] = 64'h000000002eec1a7b;
assign WBL_ROM8[4] = 64'h000000001c5f1bf2;
assign WBL_ROM8[5] = 64'h00000000a6976e6b;
assign WBL_ROM8[6] = 64'h00000000b4445a6f;
assign WBL_ROM8[7] = 64'h00000000c617a0c5;
assign WBL_ROM8[8] = 64'h00000000e8c45230;
assign WBL_ROM8[9] = 64'h00000000dda73b01;
assign WBL_ROM8[10] = 64'h00000000747ed667;
assign WBL_ROM8[11] = 64'h000000001f3db32b;
assign WBL_ROM8[12] = 64'h000000004b6429fe;
assign WBL_ROM8[13] = 64'h00000000bd5de3d7;
assign WBL_ROM8[14] = 64'h000000008b192fab;
assign WBL_ROM8[15] = 64'h000000008a738476;
assign WBL_ROM8[16] = 64'h00000000706053ca;
assign WBL_ROM8[17] = 64'h000000003e81d182;
assign WBL_ROM8[18] = 64'h00000000b54f00c9;
assign WBL_ROM8[19] = 64'h0000000066dced7d;
assign WBL_ROM8[20] = 64'h00000000482220fa;
assign WBL_ROM8[21] = 64'h00000000032afc59;
assign WBL_ROM8[22] = 64'h00000000f690b147;
assign WBL_ROM8[23] = 64'h000000000e885bf0;
assign WBL_ROM8[24] = 64'h0000000061466aad;
assign WBL_ROM8[25] = 64'h0000000035eecbd4;
assign WBL_ROM8[26] = 64'h0000000057b8bea2;
assign WBL_ROM8[27] = 64'h00000000b91439af;
assign WBL_ROM8[28] = 64'h0000000086de4a9c;
assign WBL_ROM8[29] = 64'h00000000c15e4ca4;
assign WBL_ROM8[30] = 64'h000000001d0b5872;
assign WBL_ROM8[31] = 64'h000000009edbcfc0;
assign WBL_ROM8[32] = 64'hff55224ee1e0d0b7;
assign WBL_ROM8[33] = 64'h9489c7caf832effd;
assign WBL_ROM8[34] = 64'h91d8d300983aaa93;
assign WBL_ROM8[35] = 64'h00000000110afb26;
assign WBL_ROM8[36] = 64'h0000000069494336;
assign WBL_ROM8[37] = 64'h00000000d9064d3f;
assign WBL_ROM8[38] = 64'h000000008e2433f7;
assign WBL_ROM8[39] = 64'h00000000945c85cc;
assign WBL_ROM8[40] = 64'h000000009bc24534;
assign WBL_ROM8[41] = 64'h000000001ed3f9a5;
assign WBL_ROM8[42] = 64'h0000000087ac02e5;
assign WBL_ROM8[43] = 64'h00000000e9627ff1;
assign WBL_ROM8[44] = 64'h00000000ce915071;
assign WBL_ROM8[45] = 64'h0000000055953cd8;
assign WBL_ROM8[46] = 64'h0000000028e49f31;
assign WBL_ROM8[47] = 64'h00000000df79a815;
assign WBL_ROM8[48] = 64'h000000008ce75104;
assign WBL_ROM8[49] = 64'h00000000a1c8a3c7;
assign WBL_ROM8[50] = 64'h0000000089374023;
assign WBL_ROM8[51] = 64'h000000000d6d8fc3;
assign WBL_ROM8[52] = 64'h00000000bf8d9218;
assign WBL_ROM8[53] = 64'h00000000e6d59d96;
assign WBL_ROM8[54] = 64'h00000000424e3805;
assign WBL_ROM8[55] = 64'h0000000068a9f59a;
assign WBL_ROM8[56] = 64'h00000000416cbc07;
assign WBL_ROM8[57] = 64'h000000009956b612;
assign WBL_ROM8[58] = 64'h000000002df4da80;
assign WBL_ROM8[59] = 64'h000000000fea21e2;
assign WBL_ROM8[60] = 64'h00000000b06510eb;
assign WBL_ROM8[61] = 64'h00000000547aff27;
assign WBL_ROM8[62] = 64'h00000000bbaef3b2;
assign WBL_ROM8[63] = 64'h000000001608d275;

wire [63:0] WBL_ROM9 [0:63];
assign WBL_ROM9[0] = 64'hff66789fbacd0963;
assign WBL_ROM9[1] = 64'hb33ccfa6780c837c;
assign WBL_ROM9[2] = 64'hd2e8df0025132c77;
assign WBL_ROM9[3] = 64'h000000002eec1a7b;
assign WBL_ROM9[4] = 64'h000000001c5f1bf2;
assign WBL_ROM9[5] = 64'h00000000a6976e6b;
assign WBL_ROM9[6] = 64'h00000000b4445a6f;
assign WBL_ROM9[7] = 64'h00000000c617a0c5;
assign WBL_ROM9[8] = 64'h00000000e8c45230;
assign WBL_ROM9[9] = 64'h00000000dda73b01;
assign WBL_ROM9[10] = 64'h00000000747ed667;
assign WBL_ROM9[11] = 64'h000000001f3db32b;
assign WBL_ROM9[12] = 64'h000000004b6429fe;
assign WBL_ROM9[13] = 64'h00000000bd5de3d7;
assign WBL_ROM9[14] = 64'h000000008b192fab;
assign WBL_ROM9[15] = 64'h000000008a738476;
assign WBL_ROM9[16] = 64'h00000000706053ca;
assign WBL_ROM9[17] = 64'h000000003e81d182;
assign WBL_ROM9[18] = 64'h00000000b54f00c9;
assign WBL_ROM9[19] = 64'h0000000066dced7d;
assign WBL_ROM9[20] = 64'h00000000482220fa;
assign WBL_ROM9[21] = 64'h00000000032afc59;
assign WBL_ROM9[22] = 64'h00000000f690b147;
assign WBL_ROM9[23] = 64'h000000000e885bf0;
assign WBL_ROM9[24] = 64'h0000000061466aad;
assign WBL_ROM9[25] = 64'h0000000035eecbd4;
assign WBL_ROM9[26] = 64'h0000000057b8bea2;
assign WBL_ROM9[27] = 64'h00000000b91439af;
assign WBL_ROM9[28] = 64'h0000000086de4a9c;
assign WBL_ROM9[29] = 64'h00000000c15e4ca4;
assign WBL_ROM9[30] = 64'h000000001d0b5872;
assign WBL_ROM9[31] = 64'h000000009edbcfc0;
assign WBL_ROM9[32] = 64'h00998760e1e0d0b7;
assign WBL_ROM9[33] = 64'h4cc33059f832effd;
assign WBL_ROM9[34] = 64'h2d172000983aaa93;
assign WBL_ROM9[35] = 64'h00000000110afb26;
assign WBL_ROM9[36] = 64'h0000000069494336;
assign WBL_ROM9[37] = 64'h00000000d9064d3f;
assign WBL_ROM9[38] = 64'h000000008e2433f7;
assign WBL_ROM9[39] = 64'h00000000945c85cc;
assign WBL_ROM9[40] = 64'h000000009bc24534;
assign WBL_ROM9[41] = 64'h000000001ed3f9a5;
assign WBL_ROM9[42] = 64'h0000000087ac02e5;
assign WBL_ROM9[43] = 64'h00000000e9627ff1;
assign WBL_ROM9[44] = 64'h00000000ce915071;
assign WBL_ROM9[45] = 64'h0000000055953cd8;
assign WBL_ROM9[46] = 64'h0000000028e49f31;
assign WBL_ROM9[47] = 64'h00000000df79a815;
assign WBL_ROM9[48] = 64'h000000008ce75104;
assign WBL_ROM9[49] = 64'h00000000a1c8a3c7;
assign WBL_ROM9[50] = 64'h0000000089374023;
assign WBL_ROM9[51] = 64'h000000000d6d8fc3;
assign WBL_ROM9[52] = 64'h00000000bf8d9218;
assign WBL_ROM9[53] = 64'h00000000e6d59d96;
assign WBL_ROM9[54] = 64'h00000000424e3805;
assign WBL_ROM9[55] = 64'h0000000068a9f59a;
assign WBL_ROM9[56] = 64'h00000000416cbc07;
assign WBL_ROM9[57] = 64'h000000009956b612;
assign WBL_ROM9[58] = 64'h000000002df4da80;
assign WBL_ROM9[59] = 64'h000000000fea21e2;
assign WBL_ROM9[60] = 64'h00000000b06510eb;
assign WBL_ROM9[61] = 64'h00000000547aff27;
assign WBL_ROM9[62] = 64'h00000000bbaef3b2;
assign WBL_ROM9[63] = 64'h000000001608d275;

wire [63:0] WBL_ROM10 [0:63];
assign WBL_ROM10[0] = 64'h55bbc9f4bacd0963;
assign WBL_ROM10[1] = 64'h90bf3369780c837c;
assign WBL_ROM10[2] = 64'h8b095e0025132c77;
assign WBL_ROM10[3] = 64'h000000002eec1a7b;
assign WBL_ROM10[4] = 64'h000000001c5f1bf2;
assign WBL_ROM10[5] = 64'h00000000a6976e6b;
assign WBL_ROM10[6] = 64'h00000000b4445a6f;
assign WBL_ROM10[7] = 64'h00000000c617a0c5;
assign WBL_ROM10[8] = 64'h00000000e8c45230;
assign WBL_ROM10[9] = 64'h00000000dda73b01;
assign WBL_ROM10[10] = 64'h00000000747ed667;
assign WBL_ROM10[11] = 64'h000000001f3db32b;
assign WBL_ROM10[12] = 64'h000000004b6429fe;
assign WBL_ROM10[13] = 64'h00000000bd5de3d7;
assign WBL_ROM10[14] = 64'h000000008b192fab;
assign WBL_ROM10[15] = 64'h000000008a738476;
assign WBL_ROM10[16] = 64'h00000000706053ca;
assign WBL_ROM10[17] = 64'h000000003e81d182;
assign WBL_ROM10[18] = 64'h00000000b54f00c9;
assign WBL_ROM10[19] = 64'h0000000066dced7d;
assign WBL_ROM10[20] = 64'h00000000482220fa;
assign WBL_ROM10[21] = 64'h00000000032afc59;
assign WBL_ROM10[22] = 64'h00000000f690b147;
assign WBL_ROM10[23] = 64'h000000000e885bf0;
assign WBL_ROM10[24] = 64'h0000000061466aad;
assign WBL_ROM10[25] = 64'h0000000035eecbd4;
assign WBL_ROM10[26] = 64'h0000000057b8bea2;
assign WBL_ROM10[27] = 64'h00000000b91439af;
assign WBL_ROM10[28] = 64'h0000000086de4a9c;
assign WBL_ROM10[29] = 64'h00000000c15e4ca4;
assign WBL_ROM10[30] = 64'h000000001d0b5872;
assign WBL_ROM10[31] = 64'h000000009edbcfc0;
assign WBL_ROM10[32] = 64'haa44360be1e0d0b7;
assign WBL_ROM10[33] = 64'h6f40cc96f832effd;
assign WBL_ROM10[34] = 64'h74f6a100983aaa93;
assign WBL_ROM10[35] = 64'h00000000110afb26;
assign WBL_ROM10[36] = 64'h0000000069494336;
assign WBL_ROM10[37] = 64'h00000000d9064d3f;
assign WBL_ROM10[38] = 64'h000000008e2433f7;
assign WBL_ROM10[39] = 64'h00000000945c85cc;
assign WBL_ROM10[40] = 64'h000000009bc24534;
assign WBL_ROM10[41] = 64'h000000001ed3f9a5;
assign WBL_ROM10[42] = 64'h0000000087ac02e5;
assign WBL_ROM10[43] = 64'h00000000e9627ff1;
assign WBL_ROM10[44] = 64'h00000000ce915071;
assign WBL_ROM10[45] = 64'h0000000055953cd8;
assign WBL_ROM10[46] = 64'h0000000028e49f31;
assign WBL_ROM10[47] = 64'h00000000df79a815;
assign WBL_ROM10[48] = 64'h000000008ce75104;
assign WBL_ROM10[49] = 64'h00000000a1c8a3c7;
assign WBL_ROM10[50] = 64'h0000000089374023;
assign WBL_ROM10[51] = 64'h000000000d6d8fc3;
assign WBL_ROM10[52] = 64'h00000000bf8d9218;
assign WBL_ROM10[53] = 64'h00000000e6d59d96;
assign WBL_ROM10[54] = 64'h00000000424e3805;
assign WBL_ROM10[55] = 64'h0000000068a9f59a;
assign WBL_ROM10[56] = 64'h00000000416cbc07;
assign WBL_ROM10[57] = 64'h000000009956b612;
assign WBL_ROM10[58] = 64'h000000002df4da80;
assign WBL_ROM10[59] = 64'h000000000fea21e2;
assign WBL_ROM10[60] = 64'h00000000b06510eb;
assign WBL_ROM10[61] = 64'h00000000547aff27;
assign WBL_ROM10[62] = 64'h00000000bbaef3b2;
assign WBL_ROM10[63] = 64'h000000001608d275;

wire [63:0] WBL_ROM11 [0:63];
assign WBL_ROM11[0] = 64'h336921d4bacd0963;
assign WBL_ROM11[1] = 64'hef267835780c837c;
assign WBL_ROM11[2] = 64'h6e27790025132c77;
assign WBL_ROM11[3] = 64'h000000002eec1a7b;
assign WBL_ROM11[4] = 64'h000000001c5f1bf2;
assign WBL_ROM11[5] = 64'h00000000a6976e6b;
assign WBL_ROM11[6] = 64'h00000000b4445a6f;
assign WBL_ROM11[7] = 64'h00000000c617a0c5;
assign WBL_ROM11[8] = 64'h00000000e8c45230;
assign WBL_ROM11[9] = 64'h00000000dda73b01;
assign WBL_ROM11[10] = 64'h00000000747ed667;
assign WBL_ROM11[11] = 64'h000000001f3db32b;
assign WBL_ROM11[12] = 64'h000000004b6429fe;
assign WBL_ROM11[13] = 64'h00000000bd5de3d7;
assign WBL_ROM11[14] = 64'h000000008b192fab;
assign WBL_ROM11[15] = 64'h000000008a738476;
assign WBL_ROM11[16] = 64'h00000000706053ca;
assign WBL_ROM11[17] = 64'h000000003e81d182;
assign WBL_ROM11[18] = 64'h00000000b54f00c9;
assign WBL_ROM11[19] = 64'h0000000066dced7d;
assign WBL_ROM11[20] = 64'h00000000482220fa;
assign WBL_ROM11[21] = 64'h00000000032afc59;
assign WBL_ROM11[22] = 64'h00000000f690b147;
assign WBL_ROM11[23] = 64'h000000000e885bf0;
assign WBL_ROM11[24] = 64'h0000000061466aad;
assign WBL_ROM11[25] = 64'h0000000035eecbd4;
assign WBL_ROM11[26] = 64'h0000000057b8bea2;
assign WBL_ROM11[27] = 64'h00000000b91439af;
assign WBL_ROM11[28] = 64'h0000000086de4a9c;
assign WBL_ROM11[29] = 64'h00000000c15e4ca4;
assign WBL_ROM11[30] = 64'h000000001d0b5872;
assign WBL_ROM11[31] = 64'h000000009edbcfc0;
assign WBL_ROM11[32] = 64'hcc96de2be1e0d0b7;
assign WBL_ROM11[33] = 64'h10d987caf832effd;
assign WBL_ROM11[34] = 64'h91d88600983aaa93;
assign WBL_ROM11[35] = 64'h00000000110afb26;
assign WBL_ROM11[36] = 64'h0000000069494336;
assign WBL_ROM11[37] = 64'h00000000d9064d3f;
assign WBL_ROM11[38] = 64'h000000008e2433f7;
assign WBL_ROM11[39] = 64'h00000000945c85cc;
assign WBL_ROM11[40] = 64'h000000009bc24534;
assign WBL_ROM11[41] = 64'h000000001ed3f9a5;
assign WBL_ROM11[42] = 64'h0000000087ac02e5;
assign WBL_ROM11[43] = 64'h00000000e9627ff1;
assign WBL_ROM11[44] = 64'h00000000ce915071;
assign WBL_ROM11[45] = 64'h0000000055953cd8;
assign WBL_ROM11[46] = 64'h0000000028e49f31;
assign WBL_ROM11[47] = 64'h00000000df79a815;
assign WBL_ROM11[48] = 64'h000000008ce75104;
assign WBL_ROM11[49] = 64'h00000000a1c8a3c7;
assign WBL_ROM11[50] = 64'h0000000089374023;
assign WBL_ROM11[51] = 64'h000000000d6d8fc3;
assign WBL_ROM11[52] = 64'h00000000bf8d9218;
assign WBL_ROM11[53] = 64'h00000000e6d59d96;
assign WBL_ROM11[54] = 64'h00000000424e3805;
assign WBL_ROM11[55] = 64'h0000000068a9f59a;
assign WBL_ROM11[56] = 64'h00000000416cbc07;
assign WBL_ROM11[57] = 64'h000000009956b612;
assign WBL_ROM11[58] = 64'h000000002df4da80;
assign WBL_ROM11[59] = 64'h000000000fea21e2;
assign WBL_ROM11[60] = 64'h00000000b06510eb;
assign WBL_ROM11[61] = 64'h00000000547aff27;
assign WBL_ROM11[62] = 64'h00000000bbaef3b2;
assign WBL_ROM11[63] = 64'h000000001608d275;

wire [63:0] WBL_ROM12 [0:63];
assign WBL_ROM12[0] = 64'h0ff369debacd0963;
assign WBL_ROM12[1] = 64'h4df1c1fe780c837c;
assign WBL_ROM12[2] = 64'h3297460025132c77;
assign WBL_ROM12[3] = 64'h000000002eec1a7b;
assign WBL_ROM12[4] = 64'h000000001c5f1bf2;
assign WBL_ROM12[5] = 64'h00000000a6976e6b;
assign WBL_ROM12[6] = 64'h00000000b4445a6f;
assign WBL_ROM12[7] = 64'h00000000c617a0c5;
assign WBL_ROM12[8] = 64'h00000000e8c45230;
assign WBL_ROM12[9] = 64'h00000000dda73b01;
assign WBL_ROM12[10] = 64'h00000000747ed667;
assign WBL_ROM12[11] = 64'h000000001f3db32b;
assign WBL_ROM12[12] = 64'h000000004b6429fe;
assign WBL_ROM12[13] = 64'h00000000bd5de3d7;
assign WBL_ROM12[14] = 64'h000000008b192fab;
assign WBL_ROM12[15] = 64'h000000008a738476;
assign WBL_ROM12[16] = 64'h00000000706053ca;
assign WBL_ROM12[17] = 64'h000000003e81d182;
assign WBL_ROM12[18] = 64'h00000000b54f00c9;
assign WBL_ROM12[19] = 64'h0000000066dced7d;
assign WBL_ROM12[20] = 64'h00000000482220fa;
assign WBL_ROM12[21] = 64'h00000000032afc59;
assign WBL_ROM12[22] = 64'h00000000f690b147;
assign WBL_ROM12[23] = 64'h000000000e885bf0;
assign WBL_ROM12[24] = 64'h0000000061466aad;
assign WBL_ROM12[25] = 64'h0000000035eecbd4;
assign WBL_ROM12[26] = 64'h0000000057b8bea2;
assign WBL_ROM12[27] = 64'h00000000b91439af;
assign WBL_ROM12[28] = 64'h0000000086de4a9c;
assign WBL_ROM12[29] = 64'h00000000c15e4ca4;
assign WBL_ROM12[30] = 64'h000000001d0b5872;
assign WBL_ROM12[31] = 64'h000000009edbcfc0;
assign WBL_ROM12[32] = 64'hf00c9621e1e0d0b7;
assign WBL_ROM12[33] = 64'hb20e3e01f832effd;
assign WBL_ROM12[34] = 64'hcd68b900983aaa93;
assign WBL_ROM12[35] = 64'h00000000110afb26;
assign WBL_ROM12[36] = 64'h0000000069494336;
assign WBL_ROM12[37] = 64'h00000000d9064d3f;
assign WBL_ROM12[38] = 64'h000000008e2433f7;
assign WBL_ROM12[39] = 64'h00000000945c85cc;
assign WBL_ROM12[40] = 64'h000000009bc24534;
assign WBL_ROM12[41] = 64'h000000001ed3f9a5;
assign WBL_ROM12[42] = 64'h0000000087ac02e5;
assign WBL_ROM12[43] = 64'h00000000e9627ff1;
assign WBL_ROM12[44] = 64'h00000000ce915071;
assign WBL_ROM12[45] = 64'h0000000055953cd8;
assign WBL_ROM12[46] = 64'h0000000028e49f31;
assign WBL_ROM12[47] = 64'h00000000df79a815;
assign WBL_ROM12[48] = 64'h000000008ce75104;
assign WBL_ROM12[49] = 64'h00000000a1c8a3c7;
assign WBL_ROM12[50] = 64'h0000000089374023;
assign WBL_ROM12[51] = 64'h000000000d6d8fc3;
assign WBL_ROM12[52] = 64'h00000000bf8d9218;
assign WBL_ROM12[53] = 64'h00000000e6d59d96;
assign WBL_ROM12[54] = 64'h00000000424e3805;
assign WBL_ROM12[55] = 64'h0000000068a9f59a;
assign WBL_ROM12[56] = 64'h00000000416cbc07;
assign WBL_ROM12[57] = 64'h000000009956b612;
assign WBL_ROM12[58] = 64'h000000002df4da80;
assign WBL_ROM12[59] = 64'h000000000fea21e2;
assign WBL_ROM12[60] = 64'h00000000b06510eb;
assign WBL_ROM12[61] = 64'h00000000547aff27;
assign WBL_ROM12[62] = 64'h00000000bbaef3b2;
assign WBL_ROM12[63] = 64'h000000001608d275;

wire [63:0] WBL_ROM13 [0:63];
assign WBL_ROM13[0] = 64'h0055bb9cbacd0963;
assign WBL_ROM13[1] = 64'he52ed8e0780c837c;
assign WBL_ROM13[2] = 64'h7fccf00025132c77;
assign WBL_ROM13[3] = 64'h000000002eec1a7b;
assign WBL_ROM13[4] = 64'h000000001c5f1bf2;
assign WBL_ROM13[5] = 64'h00000000a6976e6b;
assign WBL_ROM13[6] = 64'h00000000b4445a6f;
assign WBL_ROM13[7] = 64'h00000000c617a0c5;
assign WBL_ROM13[8] = 64'h00000000e8c45230;
assign WBL_ROM13[9] = 64'h00000000dda73b01;
assign WBL_ROM13[10] = 64'h00000000747ed667;
assign WBL_ROM13[11] = 64'h000000001f3db32b;
assign WBL_ROM13[12] = 64'h000000004b6429fe;
assign WBL_ROM13[13] = 64'h00000000bd5de3d7;
assign WBL_ROM13[14] = 64'h000000008b192fab;
assign WBL_ROM13[15] = 64'h000000008a738476;
assign WBL_ROM13[16] = 64'h00000000706053ca;
assign WBL_ROM13[17] = 64'h000000003e81d182;
assign WBL_ROM13[18] = 64'h00000000b54f00c9;
assign WBL_ROM13[19] = 64'h0000000066dced7d;
assign WBL_ROM13[20] = 64'h00000000482220fa;
assign WBL_ROM13[21] = 64'h00000000032afc59;
assign WBL_ROM13[22] = 64'h00000000f690b147;
assign WBL_ROM13[23] = 64'h000000000e885bf0;
assign WBL_ROM13[24] = 64'h0000000061466aad;
assign WBL_ROM13[25] = 64'h0000000035eecbd4;
assign WBL_ROM13[26] = 64'h0000000057b8bea2;
assign WBL_ROM13[27] = 64'h00000000b91439af;
assign WBL_ROM13[28] = 64'h0000000086de4a9c;
assign WBL_ROM13[29] = 64'h00000000c15e4ca4;
assign WBL_ROM13[30] = 64'h000000001d0b5872;
assign WBL_ROM13[31] = 64'h000000009edbcfc0;
assign WBL_ROM13[32] = 64'hffaa4463e1e0d0b7;
assign WBL_ROM13[33] = 64'h1ad1271ff832effd;
assign WBL_ROM13[34] = 64'h80330f00983aaa93;
assign WBL_ROM13[35] = 64'h00000000110afb26;
assign WBL_ROM13[36] = 64'h0000000069494336;
assign WBL_ROM13[37] = 64'h00000000d9064d3f;
assign WBL_ROM13[38] = 64'h000000008e2433f7;
assign WBL_ROM13[39] = 64'h00000000945c85cc;
assign WBL_ROM13[40] = 64'h000000009bc24534;
assign WBL_ROM13[41] = 64'h000000001ed3f9a5;
assign WBL_ROM13[42] = 64'h0000000087ac02e5;
assign WBL_ROM13[43] = 64'h00000000e9627ff1;
assign WBL_ROM13[44] = 64'h00000000ce915071;
assign WBL_ROM13[45] = 64'h0000000055953cd8;
assign WBL_ROM13[46] = 64'h0000000028e49f31;
assign WBL_ROM13[47] = 64'h00000000df79a815;
assign WBL_ROM13[48] = 64'h000000008ce75104;
assign WBL_ROM13[49] = 64'h00000000a1c8a3c7;
assign WBL_ROM13[50] = 64'h0000000089374023;
assign WBL_ROM13[51] = 64'h000000000d6d8fc3;
assign WBL_ROM13[52] = 64'h00000000bf8d9218;
assign WBL_ROM13[53] = 64'h00000000e6d59d96;
assign WBL_ROM13[54] = 64'h00000000424e3805;
assign WBL_ROM13[55] = 64'h0000000068a9f59a;
assign WBL_ROM13[56] = 64'h00000000416cbc07;
assign WBL_ROM13[57] = 64'h000000009956b612;
assign WBL_ROM13[58] = 64'h000000002df4da80;
assign WBL_ROM13[59] = 64'h000000000fea21e2;
assign WBL_ROM13[60] = 64'h00000000b06510eb;
assign WBL_ROM13[61] = 64'h00000000547aff27;
assign WBL_ROM13[62] = 64'h00000000bbaef3b2;
assign WBL_ROM13[63] = 64'h000000001608d275;

wire [63:0] WBL_ROM14 [0:63];
assign WBL_ROM14[0] = 64'h00ff3396bacd0963;
assign WBL_ROM14[1] = 64'heddbe383780c837c;
assign WBL_ROM14[2] = 64'h5612420025132c77;
assign WBL_ROM14[3] = 64'h000000002eec1a7b;
assign WBL_ROM14[4] = 64'h000000001c5f1bf2;
assign WBL_ROM14[5] = 64'h00000000a6976e6b;
assign WBL_ROM14[6] = 64'h00000000b4445a6f;
assign WBL_ROM14[7] = 64'h00000000c617a0c5;
assign WBL_ROM14[8] = 64'h00000000e8c45230;
assign WBL_ROM14[9] = 64'h00000000dda73b01;
assign WBL_ROM14[10] = 64'h00000000747ed667;
assign WBL_ROM14[11] = 64'h000000001f3db32b;
assign WBL_ROM14[12] = 64'h000000004b6429fe;
assign WBL_ROM14[13] = 64'h00000000bd5de3d7;
assign WBL_ROM14[14] = 64'h000000008b192fab;
assign WBL_ROM14[15] = 64'h000000008a738476;
assign WBL_ROM14[16] = 64'h00000000706053ca;
assign WBL_ROM14[17] = 64'h000000003e81d182;
assign WBL_ROM14[18] = 64'h00000000b54f00c9;
assign WBL_ROM14[19] = 64'h0000000066dced7d;
assign WBL_ROM14[20] = 64'h00000000482220fa;
assign WBL_ROM14[21] = 64'h00000000032afc59;
assign WBL_ROM14[22] = 64'h00000000f690b147;
assign WBL_ROM14[23] = 64'h000000000e885bf0;
assign WBL_ROM14[24] = 64'h0000000061466aad;
assign WBL_ROM14[25] = 64'h0000000035eecbd4;
assign WBL_ROM14[26] = 64'h0000000057b8bea2;
assign WBL_ROM14[27] = 64'h00000000b91439af;
assign WBL_ROM14[28] = 64'h0000000086de4a9c;
assign WBL_ROM14[29] = 64'h00000000c15e4ca4;
assign WBL_ROM14[30] = 64'h000000001d0b5872;
assign WBL_ROM14[31] = 64'h000000009edbcfc0;
assign WBL_ROM14[32] = 64'hff00cc69e1e0d0b7;
assign WBL_ROM14[33] = 64'h12241c7cf832effd;
assign WBL_ROM14[34] = 64'ha9edbd00983aaa93;
assign WBL_ROM14[35] = 64'h00000000110afb26;
assign WBL_ROM14[36] = 64'h0000000069494336;
assign WBL_ROM14[37] = 64'h00000000d9064d3f;
assign WBL_ROM14[38] = 64'h000000008e2433f7;
assign WBL_ROM14[39] = 64'h00000000945c85cc;
assign WBL_ROM14[40] = 64'h000000009bc24534;
assign WBL_ROM14[41] = 64'h000000001ed3f9a5;
assign WBL_ROM14[42] = 64'h0000000087ac02e5;
assign WBL_ROM14[43] = 64'h00000000e9627ff1;
assign WBL_ROM14[44] = 64'h00000000ce915071;
assign WBL_ROM14[45] = 64'h0000000055953cd8;
assign WBL_ROM14[46] = 64'h0000000028e49f31;
assign WBL_ROM14[47] = 64'h00000000df79a815;
assign WBL_ROM14[48] = 64'h000000008ce75104;
assign WBL_ROM14[49] = 64'h00000000a1c8a3c7;
assign WBL_ROM14[50] = 64'h0000000089374023;
assign WBL_ROM14[51] = 64'h000000000d6d8fc3;
assign WBL_ROM14[52] = 64'h00000000bf8d9218;
assign WBL_ROM14[53] = 64'h00000000e6d59d96;
assign WBL_ROM14[54] = 64'h00000000424e3805;
assign WBL_ROM14[55] = 64'h0000000068a9f59a;
assign WBL_ROM14[56] = 64'h00000000416cbc07;
assign WBL_ROM14[57] = 64'h000000009956b612;
assign WBL_ROM14[58] = 64'h000000002df4da80;
assign WBL_ROM14[59] = 64'h000000000fea21e2;
assign WBL_ROM14[60] = 64'h00000000b06510eb;
assign WBL_ROM14[61] = 64'h00000000547aff27;
assign WBL_ROM14[62] = 64'h00000000bbaef3b2;
assign WBL_ROM14[63] = 64'h000000001608d275;

wire [63:0] WBL_ROM15 [0:63];
assign WBL_ROM15[0] = 64'h005511ebbacd0963;
assign WBL_ROM15[1] = 64'h895e4da4780c837c;
assign WBL_ROM15[2] = 64'h8551410025132c77;
assign WBL_ROM15[3] = 64'h000000002eec1a7b;
assign WBL_ROM15[4] = 64'h000000001c5f1bf2;
assign WBL_ROM15[5] = 64'h00000000a6976e6b;
assign WBL_ROM15[6] = 64'h00000000b4445a6f;
assign WBL_ROM15[7] = 64'h00000000c617a0c5;
assign WBL_ROM15[8] = 64'h00000000e8c45230;
assign WBL_ROM15[9] = 64'h00000000dda73b01;
assign WBL_ROM15[10] = 64'h00000000747ed667;
assign WBL_ROM15[11] = 64'h000000001f3db32b;
assign WBL_ROM15[12] = 64'h000000004b6429fe;
assign WBL_ROM15[13] = 64'h00000000bd5de3d7;
assign WBL_ROM15[14] = 64'h000000008b192fab;
assign WBL_ROM15[15] = 64'h000000008a738476;
assign WBL_ROM15[16] = 64'h00000000706053ca;
assign WBL_ROM15[17] = 64'h000000003e81d182;
assign WBL_ROM15[18] = 64'h00000000b54f00c9;
assign WBL_ROM15[19] = 64'h0000000066dced7d;
assign WBL_ROM15[20] = 64'h00000000482220fa;
assign WBL_ROM15[21] = 64'h00000000032afc59;
assign WBL_ROM15[22] = 64'h00000000f690b147;
assign WBL_ROM15[23] = 64'h000000000e885bf0;
assign WBL_ROM15[24] = 64'h0000000061466aad;
assign WBL_ROM15[25] = 64'h0000000035eecbd4;
assign WBL_ROM15[26] = 64'h0000000057b8bea2;
assign WBL_ROM15[27] = 64'h00000000b91439af;
assign WBL_ROM15[28] = 64'h0000000086de4a9c;
assign WBL_ROM15[29] = 64'h00000000c15e4ca4;
assign WBL_ROM15[30] = 64'h000000001d0b5872;
assign WBL_ROM15[31] = 64'h000000009edbcfc0;
assign WBL_ROM15[32] = 64'hffaaee14e1e0d0b7;
assign WBL_ROM15[33] = 64'h76a1b25bf832effd;
assign WBL_ROM15[34] = 64'h7aaebe00983aaa93;
assign WBL_ROM15[35] = 64'h00000000110afb26;
assign WBL_ROM15[36] = 64'h0000000069494336;
assign WBL_ROM15[37] = 64'h00000000d9064d3f;
assign WBL_ROM15[38] = 64'h000000008e2433f7;
assign WBL_ROM15[39] = 64'h00000000945c85cc;
assign WBL_ROM15[40] = 64'h000000009bc24534;
assign WBL_ROM15[41] = 64'h000000001ed3f9a5;
assign WBL_ROM15[42] = 64'h0000000087ac02e5;
assign WBL_ROM15[43] = 64'h00000000e9627ff1;
assign WBL_ROM15[44] = 64'h00000000ce915071;
assign WBL_ROM15[45] = 64'h0000000055953cd8;
assign WBL_ROM15[46] = 64'h0000000028e49f31;
assign WBL_ROM15[47] = 64'h00000000df79a815;
assign WBL_ROM15[48] = 64'h000000008ce75104;
assign WBL_ROM15[49] = 64'h00000000a1c8a3c7;
assign WBL_ROM15[50] = 64'h0000000089374023;
assign WBL_ROM15[51] = 64'h000000000d6d8fc3;
assign WBL_ROM15[52] = 64'h00000000bf8d9218;
assign WBL_ROM15[53] = 64'h00000000e6d59d96;
assign WBL_ROM15[54] = 64'h00000000424e3805;
assign WBL_ROM15[55] = 64'h0000000068a9f59a;
assign WBL_ROM15[56] = 64'h00000000416cbc07;
assign WBL_ROM15[57] = 64'h000000009956b612;
assign WBL_ROM15[58] = 64'h000000002df4da80;
assign WBL_ROM15[59] = 64'h000000000fea21e2;
assign WBL_ROM15[60] = 64'h00000000b06510eb;
assign WBL_ROM15[61] = 64'h00000000547aff27;
assign WBL_ROM15[62] = 64'h00000000bbaef3b2;
assign WBL_ROM15[63] = 64'h000000001608d275;

wire [63:0] WBL_ROM16 [0:63];
assign WBL_ROM16[0] = 64'h00ff99b4bacd0963;
assign WBL_ROM16[1] = 64'hc5fb3692780c837c;
assign WBL_ROM16[2] = 64'h17ec250025132c77;
assign WBL_ROM16[3] = 64'h000000002eec1a7b;
assign WBL_ROM16[4] = 64'h000000001c5f1bf2;
assign WBL_ROM16[5] = 64'h00000000a6976e6b;
assign WBL_ROM16[6] = 64'h00000000b4445a6f;
assign WBL_ROM16[7] = 64'h00000000c617a0c5;
assign WBL_ROM16[8] = 64'h00000000e8c45230;
assign WBL_ROM16[9] = 64'h00000000dda73b01;
assign WBL_ROM16[10] = 64'h00000000747ed667;
assign WBL_ROM16[11] = 64'h000000001f3db32b;
assign WBL_ROM16[12] = 64'h000000004b6429fe;
assign WBL_ROM16[13] = 64'h00000000bd5de3d7;
assign WBL_ROM16[14] = 64'h000000008b192fab;
assign WBL_ROM16[15] = 64'h000000008a738476;
assign WBL_ROM16[16] = 64'h00000000706053ca;
assign WBL_ROM16[17] = 64'h000000003e81d182;
assign WBL_ROM16[18] = 64'h00000000b54f00c9;
assign WBL_ROM16[19] = 64'h0000000066dced7d;
assign WBL_ROM16[20] = 64'h00000000482220fa;
assign WBL_ROM16[21] = 64'h00000000032afc59;
assign WBL_ROM16[22] = 64'h00000000f690b147;
assign WBL_ROM16[23] = 64'h000000000e885bf0;
assign WBL_ROM16[24] = 64'h0000000061466aad;
assign WBL_ROM16[25] = 64'h0000000035eecbd4;
assign WBL_ROM16[26] = 64'h0000000057b8bea2;
assign WBL_ROM16[27] = 64'h00000000b91439af;
assign WBL_ROM16[28] = 64'h0000000086de4a9c;
assign WBL_ROM16[29] = 64'h00000000c15e4ca4;
assign WBL_ROM16[30] = 64'h000000001d0b5872;
assign WBL_ROM16[31] = 64'h000000009edbcfc0;
assign WBL_ROM16[32] = 64'hff00664be1e0d0b7;
assign WBL_ROM16[33] = 64'h3a04c96df832effd;
assign WBL_ROM16[34] = 64'he813da00983aaa93;
assign WBL_ROM16[35] = 64'h00000000110afb26;
assign WBL_ROM16[36] = 64'h0000000069494336;
assign WBL_ROM16[37] = 64'h00000000d9064d3f;
assign WBL_ROM16[38] = 64'h000000008e2433f7;
assign WBL_ROM16[39] = 64'h00000000945c85cc;
assign WBL_ROM16[40] = 64'h000000009bc24534;
assign WBL_ROM16[41] = 64'h000000001ed3f9a5;
assign WBL_ROM16[42] = 64'h0000000087ac02e5;
assign WBL_ROM16[43] = 64'h00000000e9627ff1;
assign WBL_ROM16[44] = 64'h00000000ce915071;
assign WBL_ROM16[45] = 64'h0000000055953cd8;
assign WBL_ROM16[46] = 64'h0000000028e49f31;
assign WBL_ROM16[47] = 64'h00000000df79a815;
assign WBL_ROM16[48] = 64'h000000008ce75104;
assign WBL_ROM16[49] = 64'h00000000a1c8a3c7;
assign WBL_ROM16[50] = 64'h0000000089374023;
assign WBL_ROM16[51] = 64'h000000000d6d8fc3;
assign WBL_ROM16[52] = 64'h00000000bf8d9218;
assign WBL_ROM16[53] = 64'h00000000e6d59d96;
assign WBL_ROM16[54] = 64'h00000000424e3805;
assign WBL_ROM16[55] = 64'h0000000068a9f59a;
assign WBL_ROM16[56] = 64'h00000000416cbc07;
assign WBL_ROM16[57] = 64'h000000009956b612;
assign WBL_ROM16[58] = 64'h000000002df4da80;
assign WBL_ROM16[59] = 64'h000000000fea21e2;
assign WBL_ROM16[60] = 64'h00000000b06510eb;
assign WBL_ROM16[61] = 64'h00000000547aff27;
assign WBL_ROM16[62] = 64'h00000000bbaef3b2;
assign WBL_ROM16[63] = 64'h000000001608d275;

